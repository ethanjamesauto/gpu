module ram
#(
    parameter Bits = 8,
    parameter AddrBits = 16
)
(
  input [(AddrBits-1):0] A,
  input [(Bits-1):0] Din,
  input str,
  input C,
  input ld,
  output [(Bits-1):0] D
);
  reg [(Bits-1):0] memory[0:((1 << AddrBits) - 1)];

  assign D = ld? memory[A] : 'hz;

  always @ (posedge C) begin
    if (str)
      memory[A] <= Din;
  end
endmodule

module rom (
    input [15:0] A,
    input sel,
    output reg [7:0] D
);
    reg [7:0] my_rom [0:6552];

    always @ (*) begin
        if (~sel)
            D = 8'hz;
        else if (A > 16'h1998)
            D = 8'h0;
        else
            D = my_rom[A];
    end

    initial begin
        my_rom[0] = 8'hc;
        my_rom[1] = 8'h0;
        my_rom[2] = 8'hff;
        my_rom[3] = 8'h0;
        my_rom[4] = 8'h0;
        my_rom[5] = 8'h41;
        my_rom[6] = 8'h0;
        my_rom[7] = 8'h0;
        my_rom[8] = 8'h0;
        my_rom[9] = 8'h0;
        my_rom[10] = 8'hff;
        my_rom[11] = 8'h0;
        my_rom[12] = 8'h0;
        my_rom[13] = 8'h40;
        my_rom[14] = 8'h0;
        my_rom[15] = 8'h0;
        my_rom[16] = 8'h0;
        my_rom[17] = 8'h50;
        my_rom[18] = 8'h8b;
        my_rom[19] = 8'h2d;
        my_rom[20] = 8'h6;
        my_rom[21] = 8'h60;
        my_rom[22] = 8'h0;
        my_rom[23] = 8'h0;
        my_rom[24] = 8'h0;
        my_rom[25] = 8'h32;
        my_rom[26] = 8'h50;
        my_rom[27] = 8'h14;
        my_rom[28] = 8'h0;
        my_rom[29] = 8'h50;
        my_rom[30] = 8'h0;
        my_rom[31] = 8'h0;
        my_rom[32] = 8'h0;
        my_rom[33] = 8'h1e;
        my_rom[34] = 8'h3c;
        my_rom[35] = 8'h30;
        my_rom[36] = 8'h0;
        my_rom[37] = 8'h50;
        my_rom[38] = 8'h0;
        my_rom[39] = 8'h0;
        my_rom[40] = 8'h1;
        my_rom[41] = 8'h0;
        my_rom[42] = 8'h0;
        my_rom[43] = 8'h0;
        my_rom[44] = 8'h0;
        my_rom[45] = 8'h0;
        my_rom[46] = 8'h0;
        my_rom[47] = 8'h0;
        my_rom[48] = 8'h0;
        my_rom[49] = 8'h0;
        my_rom[50] = 8'h0;
        my_rom[51] = 8'h0;
        my_rom[52] = 8'h0;
        my_rom[53] = 8'h0;
        my_rom[54] = 8'h0;
        my_rom[55] = 8'h0;
        my_rom[56] = 8'h0;
        my_rom[57] = 8'h0;
        my_rom[58] = 8'h0;
        my_rom[59] = 8'h0;
        my_rom[60] = 8'h0;
        my_rom[61] = 8'h0;
        my_rom[62] = 8'h0;
        my_rom[63] = 8'h0;
        my_rom[64] = 8'h74;
        my_rom[65] = 8'h18;
        my_rom[66] = 8'h0;
        my_rom[67] = 8'h0;
        my_rom[68] = 8'h0;
        my_rom[69] = 8'h0;
        my_rom[70] = 8'h0;
        my_rom[71] = 8'h0;
        my_rom[72] = 8'h0;
        my_rom[73] = 8'h0;
        my_rom[74] = 8'h0;
        my_rom[75] = 8'h0;
        my_rom[76] = 8'h0;
        my_rom[77] = 8'h0;
        my_rom[78] = 8'h0;
        my_rom[79] = 8'h0;
        my_rom[80] = 8'h8;
        my_rom[81] = 8'h8;
        my_rom[82] = 8'h8;
        my_rom[83] = 8'h8;
        my_rom[84] = 8'h8;
        my_rom[85] = 8'h8;
        my_rom[86] = 8'h8;
        my_rom[87] = 8'h8;
        my_rom[88] = 8'h8;
        my_rom[89] = 8'h8;
        my_rom[90] = 8'h49;
        my_rom[91] = 8'h49;
        my_rom[92] = 8'h49;
        my_rom[93] = 8'h49;
        my_rom[94] = 8'h8;
        my_rom[95] = 8'h8;
        my_rom[96] = 8'h8;
        my_rom[97] = 8'h8;
        my_rom[98] = 8'h8;
        my_rom[99] = 8'h8;
        my_rom[100] = 8'h8;
        my_rom[101] = 8'h8;
        my_rom[102] = 8'h8;
        my_rom[103] = 8'h8;
        my_rom[104] = 8'h8;
        my_rom[105] = 8'h8;
        my_rom[106] = 8'h8;
        my_rom[107] = 8'h8;
        my_rom[108] = 8'h8;
        my_rom[109] = 8'h8;
        my_rom[110] = 8'ha;
        my_rom[111] = 8'h8;
        my_rom[112] = 8'h8;
        my_rom[113] = 8'h8;
        my_rom[114] = 8'h8;
        my_rom[115] = 8'h8;
        my_rom[116] = 8'h8;
        my_rom[117] = 8'h49;
        my_rom[118] = 8'h49;
        my_rom[119] = 8'h49;
        my_rom[120] = 8'h49;
        my_rom[121] = 8'he1;
        my_rom[122] = 8'hf5;
        my_rom[123] = 8'hf5;
        my_rom[124] = 8'he1;
        my_rom[125] = 8'h49;
        my_rom[126] = 8'h8;
        my_rom[127] = 8'h8;
        my_rom[128] = 8'h8;
        my_rom[129] = 8'h8;
        my_rom[130] = 8'h8;
        my_rom[131] = 8'h8;
        my_rom[132] = 8'h8;
        my_rom[133] = 8'h8;
        my_rom[134] = 8'h8;
        my_rom[135] = 8'h8;
        my_rom[136] = 8'h8;
        my_rom[137] = 8'h8;
        my_rom[138] = 8'h8;
        my_rom[139] = 8'h8;
        my_rom[140] = 8'h8;
        my_rom[141] = 8'ha;
        my_rom[142] = 8'h8;
        my_rom[143] = 8'h8;
        my_rom[144] = 8'h8;
        my_rom[145] = 8'h8;
        my_rom[146] = 8'h8;
        my_rom[147] = 8'h8;
        my_rom[148] = 8'h8;
        my_rom[149] = 8'h49;
        my_rom[150] = 8'he1;
        my_rom[151] = 8'h9b;
        my_rom[152] = 8'h9b;
        my_rom[153] = 8'he1;
        my_rom[154] = 8'he1;
        my_rom[155] = 8'h9b;
        my_rom[156] = 8'h9b;
        my_rom[157] = 8'h49;
        my_rom[158] = 8'h49;
        my_rom[159] = 8'h8;
        my_rom[160] = 8'h8;
        my_rom[161] = 8'h8;
        my_rom[162] = 8'h8;
        my_rom[163] = 8'h8;
        my_rom[164] = 8'h8;
        my_rom[165] = 8'h8;
        my_rom[166] = 8'h8;
        my_rom[167] = 8'h8;
        my_rom[168] = 8'h8;
        my_rom[169] = 8'h8;
        my_rom[170] = 8'h8;
        my_rom[171] = 8'h8;
        my_rom[172] = 8'ha;
        my_rom[173] = 8'h8;
        my_rom[174] = 8'h8;
        my_rom[175] = 8'h8;
        my_rom[176] = 8'h8;
        my_rom[177] = 8'h8;
        my_rom[178] = 8'h8;
        my_rom[179] = 8'h49;
        my_rom[180] = 8'he1;
        my_rom[181] = 8'he1;
        my_rom[182] = 8'he1;
        my_rom[183] = 8'h9b;
        my_rom[184] = 8'h9b;
        my_rom[185] = 8'h9b;
        my_rom[186] = 8'h9b;
        my_rom[187] = 8'he1;
        my_rom[188] = 8'h9b;
        my_rom[189] = 8'h9b;
        my_rom[190] = 8'h49;
        my_rom[191] = 8'h8;
        my_rom[192] = 8'h8;
        my_rom[193] = 8'h8;
        my_rom[194] = 8'h8;
        my_rom[195] = 8'h8;
        my_rom[196] = 8'h8;
        my_rom[197] = 8'h8;
        my_rom[198] = 8'h8;
        my_rom[199] = 8'h8;
        my_rom[200] = 8'h8;
        my_rom[201] = 8'h8;
        my_rom[202] = 8'h8;
        my_rom[203] = 8'ha;
        my_rom[204] = 8'h8;
        my_rom[205] = 8'h8;
        my_rom[206] = 8'h8;
        my_rom[207] = 8'h8;
        my_rom[208] = 8'h8;
        my_rom[209] = 8'h49;
        my_rom[210] = 8'hf5;
        my_rom[211] = 8'he1;
        my_rom[212] = 8'he1;
        my_rom[213] = 8'h9b;
        my_rom[214] = 8'h9b;
        my_rom[215] = 8'h9b;
        my_rom[216] = 8'h9b;
        my_rom[217] = 8'he1;
        my_rom[218] = 8'he1;
        my_rom[219] = 8'hf5;
        my_rom[220] = 8'h9b;
        my_rom[221] = 8'h9b;
        my_rom[222] = 8'h49;
        my_rom[223] = 8'h8;
        my_rom[224] = 8'h8;
        my_rom[225] = 8'h8;
        my_rom[226] = 8'h8;
        my_rom[227] = 8'h8;
        my_rom[228] = 8'h8;
        my_rom[229] = 8'h8;
        my_rom[230] = 8'h8;
        my_rom[231] = 8'h8;
        my_rom[232] = 8'h8;
        my_rom[233] = 8'h8;
        my_rom[234] = 8'ha;
        my_rom[235] = 8'h8;
        my_rom[236] = 8'h8;
        my_rom[237] = 8'h8;
        my_rom[238] = 8'h8;
        my_rom[239] = 8'h49;
        my_rom[240] = 8'h9b;
        my_rom[241] = 8'hf5;
        my_rom[242] = 8'hf5;
        my_rom[243] = 8'h9b;
        my_rom[244] = 8'hf5;
        my_rom[245] = 8'he1;
        my_rom[246] = 8'hf5;
        my_rom[247] = 8'he1;
        my_rom[248] = 8'he1;
        my_rom[249] = 8'hf5;
        my_rom[250] = 8'hf5;
        my_rom[251] = 8'hf5;
        my_rom[252] = 8'h9b;
        my_rom[253] = 8'h49;
        my_rom[254] = 8'h8;
        my_rom[255] = 8'h8;
        my_rom[256] = 8'h8;
        my_rom[257] = 8'h8;
        my_rom[258] = 8'h8;
        my_rom[259] = 8'h8;
        my_rom[260] = 8'h8;
        my_rom[261] = 8'h8;
        my_rom[262] = 8'h8;
        my_rom[263] = 8'h8;
        my_rom[264] = 8'h8;
        my_rom[265] = 8'ha;
        my_rom[266] = 8'h8;
        my_rom[267] = 8'h8;
        my_rom[268] = 8'h8;
        my_rom[269] = 8'h8;
        my_rom[270] = 8'h49;
        my_rom[271] = 8'he1;
        my_rom[272] = 8'he1;
        my_rom[273] = 8'he1;
        my_rom[274] = 8'hf5;
        my_rom[275] = 8'hf5;
        my_rom[276] = 8'hf5;
        my_rom[277] = 8'hf5;
        my_rom[278] = 8'hf5;
        my_rom[279] = 8'hf5;
        my_rom[280] = 8'hf5;
        my_rom[281] = 8'he1;
        my_rom[282] = 8'he1;
        my_rom[283] = 8'h9b;
        my_rom[284] = 8'h49;
        my_rom[285] = 8'h8;
        my_rom[286] = 8'h8;
        my_rom[287] = 8'h8;
        my_rom[288] = 8'h8;
        my_rom[289] = 8'h8;
        my_rom[290] = 8'h8;
        my_rom[291] = 8'h8;
        my_rom[292] = 8'h8;
        my_rom[293] = 8'h8;
        my_rom[294] = 8'h8;
        my_rom[295] = 8'h8;
        my_rom[296] = 8'ha;
        my_rom[297] = 8'h8;
        my_rom[298] = 8'h8;
        my_rom[299] = 8'h8;
        my_rom[300] = 8'h8;
        my_rom[301] = 8'h8;
        my_rom[302] = 8'h49;
        my_rom[303] = 8'h9b;
        my_rom[304] = 8'he1;
        my_rom[305] = 8'he1;
        my_rom[306] = 8'he1;
        my_rom[307] = 8'he1;
        my_rom[308] = 8'h49;
        my_rom[309] = 8'he1;
        my_rom[310] = 8'h49;
        my_rom[311] = 8'h9b;
        my_rom[312] = 8'h9b;
        my_rom[313] = 8'he1;
        my_rom[314] = 8'h9b;
        my_rom[315] = 8'h9b;
        my_rom[316] = 8'h49;
        my_rom[317] = 8'h8;
        my_rom[318] = 8'h8;
        my_rom[319] = 8'h8;
        my_rom[320] = 8'h8;
        my_rom[321] = 8'h8;
        my_rom[322] = 8'h8;
        my_rom[323] = 8'h8;
        my_rom[324] = 8'h8;
        my_rom[325] = 8'h8;
        my_rom[326] = 8'h8;
        my_rom[327] = 8'ha;
        my_rom[328] = 8'h8;
        my_rom[329] = 8'h8;
        my_rom[330] = 8'h8;
        my_rom[331] = 8'h8;
        my_rom[332] = 8'h9b;
        my_rom[333] = 8'h49;
        my_rom[334] = 8'h9b;
        my_rom[335] = 8'he1;
        my_rom[336] = 8'he1;
        my_rom[337] = 8'h49;
        my_rom[338] = 8'h49;
        my_rom[339] = 8'heb;
        my_rom[340] = 8'h49;
        my_rom[341] = 8'heb;
        my_rom[342] = 8'h49;
        my_rom[343] = 8'h49;
        my_rom[344] = 8'h9b;
        my_rom[345] = 8'he1;
        my_rom[346] = 8'h9b;
        my_rom[347] = 8'h49;
        my_rom[348] = 8'h8;
        my_rom[349] = 8'h8;
        my_rom[350] = 8'h8;
        my_rom[351] = 8'h8;
        my_rom[352] = 8'h8;
        my_rom[353] = 8'h8;
        my_rom[354] = 8'h8;
        my_rom[355] = 8'h8;
        my_rom[356] = 8'h8;
        my_rom[357] = 8'h8;
        my_rom[358] = 8'ha;
        my_rom[359] = 8'h8;
        my_rom[360] = 8'h8;
        my_rom[361] = 8'h8;
        my_rom[362] = 8'h8;
        my_rom[363] = 8'h49;
        my_rom[364] = 8'h8;
        my_rom[365] = 8'h49;
        my_rom[366] = 8'h1;
        my_rom[367] = 8'h49;
        my_rom[368] = 8'hdb;
        my_rom[369] = 8'hdb;
        my_rom[370] = 8'hdb;
        my_rom[371] = 8'h49;
        my_rom[372] = 8'hdb;
        my_rom[373] = 8'hdb;
        my_rom[374] = 8'hdb;
        my_rom[375] = 8'h1;
        my_rom[376] = 8'h9b;
        my_rom[377] = 8'h9b;
        my_rom[378] = 8'h49;
        my_rom[379] = 8'h8;
        my_rom[380] = 8'h8;
        my_rom[381] = 8'h8;
        my_rom[382] = 8'h8;
        my_rom[383] = 8'h8;
        my_rom[384] = 8'h8;
        my_rom[385] = 8'h8;
        my_rom[386] = 8'h8;
        my_rom[387] = 8'h8;
        my_rom[388] = 8'h8;
        my_rom[389] = 8'ha;
        my_rom[390] = 8'h8;
        my_rom[391] = 8'h8;
        my_rom[392] = 8'h8;
        my_rom[393] = 8'h8;
        my_rom[394] = 8'h49;
        my_rom[395] = 8'h8;
        my_rom[396] = 8'h8;
        my_rom[397] = 8'h1;
        my_rom[398] = 8'hdb;
        my_rom[399] = 8'hff;
        my_rom[400] = 8'h1;
        my_rom[401] = 8'heb;
        my_rom[402] = 8'hdb;
        my_rom[403] = 8'h1;
        my_rom[404] = 8'hff;
        my_rom[405] = 8'hdb;
        my_rom[406] = 8'h1;
        my_rom[407] = 8'h9b;
        my_rom[408] = 8'h49;
        my_rom[409] = 8'h8;
        my_rom[410] = 8'h8;
        my_rom[411] = 8'h8;
        my_rom[412] = 8'h8;
        my_rom[413] = 8'h8;
        my_rom[414] = 8'h8;
        my_rom[415] = 8'h8;
        my_rom[416] = 8'h8;
        my_rom[417] = 8'h8;
        my_rom[418] = 8'h8;
        my_rom[419] = 8'h8;
        my_rom[420] = 8'ha;
        my_rom[421] = 8'h8;
        my_rom[422] = 8'h8;
        my_rom[423] = 8'h8;
        my_rom[424] = 8'h8;
        my_rom[425] = 8'h8;
        my_rom[426] = 8'h8;
        my_rom[427] = 8'h8;
        my_rom[428] = 8'h1;
        my_rom[429] = 8'hdb;
        my_rom[430] = 8'hff;
        my_rom[431] = 8'h1;
        my_rom[432] = 8'heb;
        my_rom[433] = 8'heb;
        my_rom[434] = 8'h1;
        my_rom[435] = 8'hff;
        my_rom[436] = 8'hdb;
        my_rom[437] = 8'h1;
        my_rom[438] = 8'h9b;
        my_rom[439] = 8'h49;
        my_rom[440] = 8'h8;
        my_rom[441] = 8'h8;
        my_rom[442] = 8'h8;
        my_rom[443] = 8'h8;
        my_rom[444] = 8'h8;
        my_rom[445] = 8'h8;
        my_rom[446] = 8'h8;
        my_rom[447] = 8'h8;
        my_rom[448] = 8'h8;
        my_rom[449] = 8'h8;
        my_rom[450] = 8'h8;
        my_rom[451] = 8'ha;
        my_rom[452] = 8'h8;
        my_rom[453] = 8'h8;
        my_rom[454] = 8'h8;
        my_rom[455] = 8'h8;
        my_rom[456] = 8'h8;
        my_rom[457] = 8'h8;
        my_rom[458] = 8'h8;
        my_rom[459] = 8'h1;
        my_rom[460] = 8'hdb;
        my_rom[461] = 8'heb;
        my_rom[462] = 8'heb;
        my_rom[463] = 8'heb;
        my_rom[464] = 8'heb;
        my_rom[465] = 8'heb;
        my_rom[466] = 8'heb;
        my_rom[467] = 8'hdb;
        my_rom[468] = 8'h1;
        my_rom[469] = 8'h49;
        my_rom[470] = 8'h8;
        my_rom[471] = 8'h8;
        my_rom[472] = 8'h8;
        my_rom[473] = 8'h8;
        my_rom[474] = 8'h8;
        my_rom[475] = 8'h8;
        my_rom[476] = 8'h8;
        my_rom[477] = 8'h8;
        my_rom[478] = 8'h8;
        my_rom[479] = 8'h8;
        my_rom[480] = 8'h8;
        my_rom[481] = 8'h8;
        my_rom[482] = 8'ha;
        my_rom[483] = 8'h8;
        my_rom[484] = 8'h8;
        my_rom[485] = 8'h8;
        my_rom[486] = 8'h8;
        my_rom[487] = 8'h8;
        my_rom[488] = 8'h8;
        my_rom[489] = 8'h45;
        my_rom[490] = 8'h45;
        my_rom[491] = 8'h1;
        my_rom[492] = 8'hdb;
        my_rom[493] = 8'heb;
        my_rom[494] = 8'heb;
        my_rom[495] = 8'heb;
        my_rom[496] = 8'heb;
        my_rom[497] = 8'hdb;
        my_rom[498] = 8'h1;
        my_rom[499] = 8'h45;
        my_rom[500] = 8'h45;
        my_rom[501] = 8'h8;
        my_rom[502] = 8'h8;
        my_rom[503] = 8'h8;
        my_rom[504] = 8'h8;
        my_rom[505] = 8'h8;
        my_rom[506] = 8'h8;
        my_rom[507] = 8'h8;
        my_rom[508] = 8'h8;
        my_rom[509] = 8'h8;
        my_rom[510] = 8'h8;
        my_rom[511] = 8'h8;
        my_rom[512] = 8'h8;
        my_rom[513] = 8'ha;
        my_rom[514] = 8'h8;
        my_rom[515] = 8'h8;
        my_rom[516] = 8'h8;
        my_rom[517] = 8'h8;
        my_rom[518] = 8'h8;
        my_rom[519] = 8'h45;
        my_rom[520] = 8'hff;
        my_rom[521] = 8'hef;
        my_rom[522] = 8'h1;
        my_rom[523] = 8'h1;
        my_rom[524] = 8'hdb;
        my_rom[525] = 8'heb;
        my_rom[526] = 8'heb;
        my_rom[527] = 8'hdb;
        my_rom[528] = 8'h1;
        my_rom[529] = 8'h1;
        my_rom[530] = 8'hff;
        my_rom[531] = 8'hef;
        my_rom[532] = 8'h45;
        my_rom[533] = 8'h8;
        my_rom[534] = 8'h8;
        my_rom[535] = 8'h8;
        my_rom[536] = 8'h8;
        my_rom[537] = 8'h8;
        my_rom[538] = 8'h8;
        my_rom[539] = 8'h8;
        my_rom[540] = 8'h8;
        my_rom[541] = 8'h8;
        my_rom[542] = 8'h8;
        my_rom[543] = 8'h8;
        my_rom[544] = 8'ha;
        my_rom[545] = 8'h8;
        my_rom[546] = 8'h8;
        my_rom[547] = 8'h8;
        my_rom[548] = 8'h8;
        my_rom[549] = 8'h8;
        my_rom[550] = 8'h45;
        my_rom[551] = 8'hef;
        my_rom[552] = 8'hef;
        my_rom[553] = 8'h9f;
        my_rom[554] = 8'h9f;
        my_rom[555] = 8'h1;
        my_rom[556] = 8'h1;
        my_rom[557] = 8'h1;
        my_rom[558] = 8'h1;
        my_rom[559] = 8'h9f;
        my_rom[560] = 8'h45;
        my_rom[561] = 8'hef;
        my_rom[562] = 8'hef;
        my_rom[563] = 8'h45;
        my_rom[564] = 8'h8;
        my_rom[565] = 8'h8;
        my_rom[566] = 8'h8;
        my_rom[567] = 8'h8;
        my_rom[568] = 8'h8;
        my_rom[569] = 8'h8;
        my_rom[570] = 8'h8;
        my_rom[571] = 8'h8;
        my_rom[572] = 8'h8;
        my_rom[573] = 8'h8;
        my_rom[574] = 8'h8;
        my_rom[575] = 8'ha;
        my_rom[576] = 8'h8;
        my_rom[577] = 8'h8;
        my_rom[578] = 8'h8;
        my_rom[579] = 8'h8;
        my_rom[580] = 8'h45;
        my_rom[581] = 8'h45;
        my_rom[582] = 8'h45;
        my_rom[583] = 8'h45;
        my_rom[584] = 8'h45;
        my_rom[585] = 8'hef;
        my_rom[586] = 8'hef;
        my_rom[587] = 8'hef;
        my_rom[588] = 8'hef;
        my_rom[589] = 8'hef;
        my_rom[590] = 8'hef;
        my_rom[591] = 8'h9f;
        my_rom[592] = 8'h45;
        my_rom[593] = 8'h45;
        my_rom[594] = 8'h45;
        my_rom[595] = 8'h45;
        my_rom[596] = 8'h8;
        my_rom[597] = 8'h8;
        my_rom[598] = 8'h8;
        my_rom[599] = 8'h8;
        my_rom[600] = 8'h8;
        my_rom[601] = 8'h8;
        my_rom[602] = 8'h8;
        my_rom[603] = 8'h8;
        my_rom[604] = 8'h8;
        my_rom[605] = 8'h8;
        my_rom[606] = 8'ha;
        my_rom[607] = 8'h8;
        my_rom[608] = 8'h8;
        my_rom[609] = 8'h8;
        my_rom[610] = 8'h8;
        my_rom[611] = 8'h45;
        my_rom[612] = 8'hdb;
        my_rom[613] = 8'hdb;
        my_rom[614] = 8'h45;
        my_rom[615] = 8'h9f;
        my_rom[616] = 8'h9f;
        my_rom[617] = 8'hef;
        my_rom[618] = 8'hff;
        my_rom[619] = 8'hff;
        my_rom[620] = 8'hff;
        my_rom[621] = 8'hef;
        my_rom[622] = 8'h9f;
        my_rom[623] = 8'h45;
        my_rom[624] = 8'h81;
        my_rom[625] = 8'hdb;
        my_rom[626] = 8'h45;
        my_rom[627] = 8'h8;
        my_rom[628] = 8'h8;
        my_rom[629] = 8'h8;
        my_rom[630] = 8'h8;
        my_rom[631] = 8'h8;
        my_rom[632] = 8'h8;
        my_rom[633] = 8'h8;
        my_rom[634] = 8'h8;
        my_rom[635] = 8'h8;
        my_rom[636] = 8'h8;
        my_rom[637] = 8'ha;
        my_rom[638] = 8'h8;
        my_rom[639] = 8'h8;
        my_rom[640] = 8'h8;
        my_rom[641] = 8'h8;
        my_rom[642] = 8'h45;
        my_rom[643] = 8'h45;
        my_rom[644] = 8'h81;
        my_rom[645] = 8'h1;
        my_rom[646] = 8'h45;
        my_rom[647] = 8'h9f;
        my_rom[648] = 8'h9f;
        my_rom[649] = 8'hef;
        my_rom[650] = 8'hef;
        my_rom[651] = 8'hef;
        my_rom[652] = 8'h9f;
        my_rom[653] = 8'h45;
        my_rom[654] = 8'h1;
        my_rom[655] = 8'h81;
        my_rom[656] = 8'h45;
        my_rom[657] = 8'h45;
        my_rom[658] = 8'h8;
        my_rom[659] = 8'h8;
        my_rom[660] = 8'h8;
        my_rom[661] = 8'h8;
        my_rom[662] = 8'h8;
        my_rom[663] = 8'h8;
        my_rom[664] = 8'h8;
        my_rom[665] = 8'h8;
        my_rom[666] = 8'h8;
        my_rom[667] = 8'h8;
        my_rom[668] = 8'ha;
        my_rom[669] = 8'h8;
        my_rom[670] = 8'h8;
        my_rom[671] = 8'h8;
        my_rom[672] = 8'h8;
        my_rom[673] = 8'h45;
        my_rom[674] = 8'h9f;
        my_rom[675] = 8'h45;
        my_rom[676] = 8'h8;
        my_rom[677] = 8'h1;
        my_rom[678] = 8'h45;
        my_rom[679] = 8'h9f;
        my_rom[680] = 8'h9f;
        my_rom[681] = 8'h9f;
        my_rom[682] = 8'h9f;
        my_rom[683] = 8'h45;
        my_rom[684] = 8'h1;
        my_rom[685] = 8'h8;
        my_rom[686] = 8'h45;
        my_rom[687] = 8'h9f;
        my_rom[688] = 8'h45;
        my_rom[689] = 8'h8;
        my_rom[690] = 8'h8;
        my_rom[691] = 8'h8;
        my_rom[692] = 8'h8;
        my_rom[693] = 8'h8;
        my_rom[694] = 8'h8;
        my_rom[695] = 8'h8;
        my_rom[696] = 8'h8;
        my_rom[697] = 8'h8;
        my_rom[698] = 8'h8;
        my_rom[699] = 8'ha;
        my_rom[700] = 8'h8;
        my_rom[701] = 8'h8;
        my_rom[702] = 8'h8;
        my_rom[703] = 8'h8;
        my_rom[704] = 8'h45;
        my_rom[705] = 8'h45;
        my_rom[706] = 8'h45;
        my_rom[707] = 8'h1;
        my_rom[708] = 8'h1;
        my_rom[709] = 8'h9f;
        my_rom[710] = 8'h45;
        my_rom[711] = 8'h45;
        my_rom[712] = 8'h45;
        my_rom[713] = 8'h45;
        my_rom[714] = 8'h9f;
        my_rom[715] = 8'h1;
        my_rom[716] = 8'h1;
        my_rom[717] = 8'h45;
        my_rom[718] = 8'h45;
        my_rom[719] = 8'h45;
        my_rom[720] = 8'h8;
        my_rom[721] = 8'h8;
        my_rom[722] = 8'h8;
        my_rom[723] = 8'h8;
        my_rom[724] = 8'h8;
        my_rom[725] = 8'h8;
        my_rom[726] = 8'h8;
        my_rom[727] = 8'h8;
        my_rom[728] = 8'h8;
        my_rom[729] = 8'h8;
        my_rom[730] = 8'ha;
        my_rom[731] = 8'h8;
        my_rom[732] = 8'h8;
        my_rom[733] = 8'h8;
        my_rom[734] = 8'h8;
        my_rom[735] = 8'h1;
        my_rom[736] = 8'heb;
        my_rom[737] = 8'heb;
        my_rom[738] = 8'h1;
        my_rom[739] = 8'h45;
        my_rom[740] = 8'h45;
        my_rom[741] = 8'h9f;
        my_rom[742] = 8'hff;
        my_rom[743] = 8'hef;
        my_rom[744] = 8'h9f;
        my_rom[745] = 8'h45;
        my_rom[746] = 8'h45;
        my_rom[747] = 8'h1;
        my_rom[748] = 8'heb;
        my_rom[749] = 8'heb;
        my_rom[750] = 8'h1;
        my_rom[751] = 8'h8;
        my_rom[752] = 8'h8;
        my_rom[753] = 8'h8;
        my_rom[754] = 8'h8;
        my_rom[755] = 8'h8;
        my_rom[756] = 8'h8;
        my_rom[757] = 8'h8;
        my_rom[758] = 8'h8;
        my_rom[759] = 8'h8;
        my_rom[760] = 8'h8;
        my_rom[761] = 8'ha;
        my_rom[762] = 8'h8;
        my_rom[763] = 8'h8;
        my_rom[764] = 8'h8;
        my_rom[765] = 8'h8;
        my_rom[766] = 8'h1;
        my_rom[767] = 8'hdb;
        my_rom[768] = 8'hdb;
        my_rom[769] = 8'h1;
        my_rom[770] = 8'h81;
        my_rom[771] = 8'h81;
        my_rom[772] = 8'h45;
        my_rom[773] = 8'h45;
        my_rom[774] = 8'h45;
        my_rom[775] = 8'h45;
        my_rom[776] = 8'h81;
        my_rom[777] = 8'h81;
        my_rom[778] = 8'h1;
        my_rom[779] = 8'hdb;
        my_rom[780] = 8'hdb;
        my_rom[781] = 8'h1;
        my_rom[782] = 8'h8;
        my_rom[783] = 8'h8;
        my_rom[784] = 8'h8;
        my_rom[785] = 8'h8;
        my_rom[786] = 8'h8;
        my_rom[787] = 8'h8;
        my_rom[788] = 8'h8;
        my_rom[789] = 8'h8;
        my_rom[790] = 8'h8;
        my_rom[791] = 8'h8;
        my_rom[792] = 8'ha;
        my_rom[793] = 8'h8;
        my_rom[794] = 8'h8;
        my_rom[795] = 8'h8;
        my_rom[796] = 8'h8;
        my_rom[797] = 8'h8;
        my_rom[798] = 8'h1;
        my_rom[799] = 8'h1;
        my_rom[800] = 8'h1;
        my_rom[801] = 8'h81;
        my_rom[802] = 8'h81;
        my_rom[803] = 8'h81;
        my_rom[804] = 8'h81;
        my_rom[805] = 8'h1;
        my_rom[806] = 8'h81;
        my_rom[807] = 8'h81;
        my_rom[808] = 8'h81;
        my_rom[809] = 8'h1;
        my_rom[810] = 8'h1;
        my_rom[811] = 8'h1;
        my_rom[812] = 8'h8;
        my_rom[813] = 8'h8;
        my_rom[814] = 8'h8;
        my_rom[815] = 8'h8;
        my_rom[816] = 8'h8;
        my_rom[817] = 8'h8;
        my_rom[818] = 8'h8;
        my_rom[819] = 8'h8;
        my_rom[820] = 8'h8;
        my_rom[821] = 8'h8;
        my_rom[822] = 8'h8;
        my_rom[823] = 8'ha;
        my_rom[824] = 8'h8;
        my_rom[825] = 8'h8;
        my_rom[826] = 8'h8;
        my_rom[827] = 8'h8;
        my_rom[828] = 8'h8;
        my_rom[829] = 8'h8;
        my_rom[830] = 8'h8;
        my_rom[831] = 8'h1;
        my_rom[832] = 8'h81;
        my_rom[833] = 8'hdb;
        my_rom[834] = 8'h81;
        my_rom[835] = 8'h81;
        my_rom[836] = 8'h1;
        my_rom[837] = 8'h81;
        my_rom[838] = 8'h81;
        my_rom[839] = 8'h81;
        my_rom[840] = 8'h1;
        my_rom[841] = 8'h8;
        my_rom[842] = 8'h8;
        my_rom[843] = 8'h8;
        my_rom[844] = 8'h8;
        my_rom[845] = 8'h8;
        my_rom[846] = 8'h8;
        my_rom[847] = 8'h8;
        my_rom[848] = 8'h8;
        my_rom[849] = 8'h8;
        my_rom[850] = 8'h8;
        my_rom[851] = 8'h8;
        my_rom[852] = 8'h8;
        my_rom[853] = 8'h8;
        my_rom[854] = 8'ha;
        my_rom[855] = 8'h8;
        my_rom[856] = 8'h8;
        my_rom[857] = 8'h8;
        my_rom[858] = 8'h8;
        my_rom[859] = 8'h8;
        my_rom[860] = 8'h8;
        my_rom[861] = 8'h8;
        my_rom[862] = 8'h1;
        my_rom[863] = 8'h81;
        my_rom[864] = 8'h81;
        my_rom[865] = 8'h81;
        my_rom[866] = 8'h81;
        my_rom[867] = 8'h1;
        my_rom[868] = 8'h81;
        my_rom[869] = 8'h81;
        my_rom[870] = 8'h81;
        my_rom[871] = 8'h1;
        my_rom[872] = 8'h8;
        my_rom[873] = 8'h8;
        my_rom[874] = 8'h8;
        my_rom[875] = 8'h8;
        my_rom[876] = 8'h8;
        my_rom[877] = 8'h8;
        my_rom[878] = 8'h8;
        my_rom[879] = 8'h8;
        my_rom[880] = 8'h8;
        my_rom[881] = 8'h8;
        my_rom[882] = 8'h8;
        my_rom[883] = 8'h8;
        my_rom[884] = 8'h8;
        my_rom[885] = 8'ha;
        my_rom[886] = 8'h8;
        my_rom[887] = 8'h8;
        my_rom[888] = 8'h8;
        my_rom[889] = 8'h8;
        my_rom[890] = 8'h8;
        my_rom[891] = 8'h8;
        my_rom[892] = 8'h8;
        my_rom[893] = 8'h8;
        my_rom[894] = 8'h1;
        my_rom[895] = 8'h81;
        my_rom[896] = 8'h81;
        my_rom[897] = 8'h81;
        my_rom[898] = 8'h1;
        my_rom[899] = 8'h81;
        my_rom[900] = 8'h81;
        my_rom[901] = 8'h1;
        my_rom[902] = 8'h8;
        my_rom[903] = 8'h8;
        my_rom[904] = 8'h8;
        my_rom[905] = 8'h8;
        my_rom[906] = 8'h8;
        my_rom[907] = 8'h8;
        my_rom[908] = 8'h8;
        my_rom[909] = 8'h8;
        my_rom[910] = 8'h8;
        my_rom[911] = 8'h8;
        my_rom[912] = 8'h8;
        my_rom[913] = 8'h8;
        my_rom[914] = 8'h8;
        my_rom[915] = 8'h8;
        my_rom[916] = 8'ha;
        my_rom[917] = 8'h8;
        my_rom[918] = 8'h8;
        my_rom[919] = 8'h8;
        my_rom[920] = 8'h8;
        my_rom[921] = 8'h8;
        my_rom[922] = 8'h8;
        my_rom[923] = 8'h8;
        my_rom[924] = 8'h8;
        my_rom[925] = 8'h1;
        my_rom[926] = 8'h81;
        my_rom[927] = 8'h81;
        my_rom[928] = 8'h81;
        my_rom[929] = 8'h1;
        my_rom[930] = 8'h81;
        my_rom[931] = 8'h81;
        my_rom[932] = 8'h1;
        my_rom[933] = 8'h8;
        my_rom[934] = 8'h8;
        my_rom[935] = 8'h8;
        my_rom[936] = 8'h8;
        my_rom[937] = 8'h8;
        my_rom[938] = 8'h8;
        my_rom[939] = 8'h8;
        my_rom[940] = 8'h8;
        my_rom[941] = 8'h8;
        my_rom[942] = 8'h8;
        my_rom[943] = 8'h8;
        my_rom[944] = 8'h8;
        my_rom[945] = 8'h8;
        my_rom[946] = 8'h8;
        my_rom[947] = 8'ha;
        my_rom[948] = 8'h8;
        my_rom[949] = 8'h8;
        my_rom[950] = 8'h8;
        my_rom[951] = 8'h8;
        my_rom[952] = 8'h8;
        my_rom[953] = 8'h8;
        my_rom[954] = 8'h8;
        my_rom[955] = 8'h8;
        my_rom[956] = 8'h1;
        my_rom[957] = 8'h9f;
        my_rom[958] = 8'h81;
        my_rom[959] = 8'h81;
        my_rom[960] = 8'h1;
        my_rom[961] = 8'h81;
        my_rom[962] = 8'h81;
        my_rom[963] = 8'h1;
        my_rom[964] = 8'h8;
        my_rom[965] = 8'h8;
        my_rom[966] = 8'h8;
        my_rom[967] = 8'h8;
        my_rom[968] = 8'h8;
        my_rom[969] = 8'h8;
        my_rom[970] = 8'h8;
        my_rom[971] = 8'h8;
        my_rom[972] = 8'h8;
        my_rom[973] = 8'h8;
        my_rom[974] = 8'h8;
        my_rom[975] = 8'h8;
        my_rom[976] = 8'h8;
        my_rom[977] = 8'h8;
        my_rom[978] = 8'ha;
        my_rom[979] = 8'h8;
        my_rom[980] = 8'h8;
        my_rom[981] = 8'h8;
        my_rom[982] = 8'h8;
        my_rom[983] = 8'h8;
        my_rom[984] = 8'h8;
        my_rom[985] = 8'h8;
        my_rom[986] = 8'h8;
        my_rom[987] = 8'h1;
        my_rom[988] = 8'hef;
        my_rom[989] = 8'hef;
        my_rom[990] = 8'h9f;
        my_rom[991] = 8'h1;
        my_rom[992] = 8'h9f;
        my_rom[993] = 8'h9f;
        my_rom[994] = 8'h1;
        my_rom[995] = 8'h8;
        my_rom[996] = 8'h8;
        my_rom[997] = 8'h8;
        my_rom[998] = 8'h8;
        my_rom[999] = 8'h8;
        my_rom[1000] = 8'h8;
        my_rom[1001] = 8'h8;
        my_rom[1002] = 8'h8;
        my_rom[1003] = 8'h8;
        my_rom[1004] = 8'h8;
        my_rom[1005] = 8'h8;
        my_rom[1006] = 8'h8;
        my_rom[1007] = 8'h8;
        my_rom[1008] = 8'h8;
        my_rom[1009] = 8'ha;
        my_rom[1010] = 8'h8;
        my_rom[1011] = 8'h8;
        my_rom[1012] = 8'h8;
        my_rom[1013] = 8'h8;
        my_rom[1014] = 8'h8;
        my_rom[1015] = 8'h8;
        my_rom[1016] = 8'h8;
        my_rom[1017] = 8'h8;
        my_rom[1018] = 8'h8;
        my_rom[1019] = 8'h1;
        my_rom[1020] = 8'h1;
        my_rom[1021] = 8'h1;
        my_rom[1022] = 8'h1;
        my_rom[1023] = 8'h1;
        my_rom[1024] = 8'h1;
        my_rom[1025] = 8'h1;
        my_rom[1026] = 8'h8;
        my_rom[1027] = 8'h8;
        my_rom[1028] = 8'h8;
        my_rom[1029] = 8'h8;
        my_rom[1030] = 8'h8;
        my_rom[1031] = 8'h8;
        my_rom[1032] = 8'h8;
        my_rom[1033] = 8'h8;
        my_rom[1034] = 8'h8;
        my_rom[1035] = 8'h8;
        my_rom[1036] = 8'h8;
        my_rom[1037] = 8'h8;
        my_rom[1038] = 8'h8;
        my_rom[1039] = 8'h8;
        my_rom[1040] = 8'ha;
        my_rom[1041] = 8'h8;
        my_rom[1042] = 8'h8;
        my_rom[1043] = 8'h8;
        my_rom[1044] = 8'h8;
        my_rom[1045] = 8'h8;
        my_rom[1046] = 8'h8;
        my_rom[1047] = 8'h8;
        my_rom[1048] = 8'h8;
        my_rom[1049] = 8'h8;
        my_rom[1050] = 8'h8;
        my_rom[1051] = 8'h8;
        my_rom[1052] = 8'h8;
        my_rom[1053] = 8'h8;
        my_rom[1054] = 8'h8;
        my_rom[1055] = 8'h8;
        my_rom[1056] = 8'h8;
        my_rom[1057] = 8'h8;
        my_rom[1058] = 8'h8;
        my_rom[1059] = 8'h8;
        my_rom[1060] = 8'h8;
        my_rom[1061] = 8'h8;
        my_rom[1062] = 8'h8;
        my_rom[1063] = 8'h8;
        my_rom[1064] = 8'h8;
        my_rom[1065] = 8'h8;
        my_rom[1066] = 8'h8;
        my_rom[1067] = 8'h8;
        my_rom[1068] = 8'h8;
        my_rom[1069] = 8'h8;
        my_rom[1070] = 8'h8;
        my_rom[1071] = 8'ha;
        my_rom[1072] = 8'h8;
        my_rom[1073] = 8'h8;
        my_rom[1074] = 8'h8;
        my_rom[1075] = 8'h8;
        my_rom[1076] = 8'h8;
        my_rom[1077] = 8'h8;
        my_rom[1078] = 8'h8;
        my_rom[1079] = 8'h8;
        my_rom[1080] = 8'h8;
        my_rom[1081] = 8'h8;
        my_rom[1082] = 8'h8;
        my_rom[1083] = 8'h8;
        my_rom[1084] = 8'h8;
        my_rom[1085] = 8'h8;
        my_rom[1086] = 8'h8;
        my_rom[1087] = 8'h8;
        my_rom[1088] = 8'h8;
        my_rom[1089] = 8'h8;
        my_rom[1090] = 8'h8;
        my_rom[1091] = 8'h8;
        my_rom[1092] = 8'h8;
        my_rom[1093] = 8'h8;
        my_rom[1094] = 8'h8;
        my_rom[1095] = 8'h8;
        my_rom[1096] = 8'h8;
        my_rom[1097] = 8'h8;
        my_rom[1098] = 8'h8;
        my_rom[1099] = 8'h8;
        my_rom[1100] = 8'h8;
        my_rom[1101] = 8'h8;
        my_rom[1102] = 8'ha;
        my_rom[1103] = 8'h8;
        my_rom[1104] = 8'h8;
        my_rom[1105] = 8'h8;
        my_rom[1106] = 8'h8;
        my_rom[1107] = 8'h8;
        my_rom[1108] = 8'h8;
        my_rom[1109] = 8'h8;
        my_rom[1110] = 8'h8;
        my_rom[1111] = 8'h8;
        my_rom[1112] = 8'h8;
        my_rom[1113] = 8'h8;
        my_rom[1114] = 8'h8;
        my_rom[1115] = 8'h8;
        my_rom[1116] = 8'h8;
        my_rom[1117] = 8'h8;
        my_rom[1118] = 8'h8;
        my_rom[1119] = 8'h8;
        my_rom[1120] = 8'h8;
        my_rom[1121] = 8'h8;
        my_rom[1122] = 8'h8;
        my_rom[1123] = 8'h8;
        my_rom[1124] = 8'h8;
        my_rom[1125] = 8'h8;
        my_rom[1126] = 8'h8;
        my_rom[1127] = 8'h8;
        my_rom[1128] = 8'h8;
        my_rom[1129] = 8'h8;
        my_rom[1130] = 8'h8;
        my_rom[1131] = 8'h8;
        my_rom[1132] = 8'h8;
        my_rom[1133] = 8'ha;
        my_rom[1134] = 8'h8;
        my_rom[1135] = 8'h8;
        my_rom[1136] = 8'h8;
        my_rom[1137] = 8'h8;
        my_rom[1138] = 8'h8;
        my_rom[1139] = 8'h8;
        my_rom[1140] = 8'h8;
        my_rom[1141] = 8'h8;
        my_rom[1142] = 8'h8;
        my_rom[1143] = 8'h8;
        my_rom[1144] = 8'h8;
        my_rom[1145] = 8'h8;
        my_rom[1146] = 8'h8;
        my_rom[1147] = 8'h8;
        my_rom[1148] = 8'h8;
        my_rom[1149] = 8'h8;
        my_rom[1150] = 8'h8;
        my_rom[1151] = 8'h8;
        my_rom[1152] = 8'h8;
        my_rom[1153] = 8'h8;
        my_rom[1154] = 8'h8;
        my_rom[1155] = 8'h8;
        my_rom[1156] = 8'h8;
        my_rom[1157] = 8'h8;
        my_rom[1158] = 8'h8;
        my_rom[1159] = 8'h8;
        my_rom[1160] = 8'h8;
        my_rom[1161] = 8'h8;
        my_rom[1162] = 8'h8;
        my_rom[1163] = 8'h8;
        my_rom[1164] = 8'ha;
        my_rom[1165] = 8'h8;
        my_rom[1166] = 8'h8;
        my_rom[1167] = 8'h8;
        my_rom[1168] = 8'h8;
        my_rom[1169] = 8'h8;
        my_rom[1170] = 8'h8;
        my_rom[1171] = 8'h8;
        my_rom[1172] = 8'h8;
        my_rom[1173] = 8'h8;
        my_rom[1174] = 8'h8;
        my_rom[1175] = 8'h8;
        my_rom[1176] = 8'h8;
        my_rom[1177] = 8'h8;
        my_rom[1178] = 8'h8;
        my_rom[1179] = 8'h8;
        my_rom[1180] = 8'h8;
        my_rom[1181] = 8'h8;
        my_rom[1182] = 8'h8;
        my_rom[1183] = 8'h8;
        my_rom[1184] = 8'h8;
        my_rom[1185] = 8'h8;
        my_rom[1186] = 8'h8;
        my_rom[1187] = 8'h8;
        my_rom[1188] = 8'h8;
        my_rom[1189] = 8'h8;
        my_rom[1190] = 8'h8;
        my_rom[1191] = 8'h8;
        my_rom[1192] = 8'h8;
        my_rom[1193] = 8'h8;
        my_rom[1194] = 8'h8;
        my_rom[1195] = 8'ha;
        my_rom[1196] = 8'h8;
        my_rom[1197] = 8'h8;
        my_rom[1198] = 8'h8;
        my_rom[1199] = 8'h8;
        my_rom[1200] = 8'h8;
        my_rom[1201] = 8'h8;
        my_rom[1202] = 8'h8;
        my_rom[1203] = 8'h8;
        my_rom[1204] = 8'h8;
        my_rom[1205] = 8'h8;
        my_rom[1206] = 8'h8;
        my_rom[1207] = 8'h8;
        my_rom[1208] = 8'h8;
        my_rom[1209] = 8'h8;
        my_rom[1210] = 8'h8;
        my_rom[1211] = 8'h8;
        my_rom[1212] = 8'h8;
        my_rom[1213] = 8'h8;
        my_rom[1214] = 8'h8;
        my_rom[1215] = 8'h8;
        my_rom[1216] = 8'h8;
        my_rom[1217] = 8'h8;
        my_rom[1218] = 8'h8;
        my_rom[1219] = 8'h8;
        my_rom[1220] = 8'h8;
        my_rom[1221] = 8'h8;
        my_rom[1222] = 8'h8;
        my_rom[1223] = 8'h8;
        my_rom[1224] = 8'h8;
        my_rom[1225] = 8'h8;
        my_rom[1226] = 8'ha;
        my_rom[1227] = 8'h8;
        my_rom[1228] = 8'h8;
        my_rom[1229] = 8'h8;
        my_rom[1230] = 8'h8;
        my_rom[1231] = 8'h8;
        my_rom[1232] = 8'h8;
        my_rom[1233] = 8'h8;
        my_rom[1234] = 8'h8;
        my_rom[1235] = 8'h8;
        my_rom[1236] = 8'h8;
        my_rom[1237] = 8'h8;
        my_rom[1238] = 8'h8;
        my_rom[1239] = 8'h8;
        my_rom[1240] = 8'h8;
        my_rom[1241] = 8'h8;
        my_rom[1242] = 8'h8;
        my_rom[1243] = 8'h8;
        my_rom[1244] = 8'h8;
        my_rom[1245] = 8'h8;
        my_rom[1246] = 8'h8;
        my_rom[1247] = 8'h8;
        my_rom[1248] = 8'h8;
        my_rom[1249] = 8'h8;
        my_rom[1250] = 8'h8;
        my_rom[1251] = 8'h8;
        my_rom[1252] = 8'h8;
        my_rom[1253] = 8'h8;
        my_rom[1254] = 8'h8;
        my_rom[1255] = 8'h8;
        my_rom[1256] = 8'h8;
        my_rom[1257] = 8'ha;
        my_rom[1258] = 8'h8;
        my_rom[1259] = 8'h8;
        my_rom[1260] = 8'h8;
        my_rom[1261] = 8'h8;
        my_rom[1262] = 8'h8;
        my_rom[1263] = 8'h8;
        my_rom[1264] = 8'h8;
        my_rom[1265] = 8'h8;
        my_rom[1266] = 8'h8;
        my_rom[1267] = 8'h8;
        my_rom[1268] = 8'h8;
        my_rom[1269] = 8'h8;
        my_rom[1270] = 8'h8;
        my_rom[1271] = 8'h8;
        my_rom[1272] = 8'h8;
        my_rom[1273] = 8'h8;
        my_rom[1274] = 8'h8;
        my_rom[1275] = 8'h8;
        my_rom[1276] = 8'h8;
        my_rom[1277] = 8'h8;
        my_rom[1278] = 8'h8;
        my_rom[1279] = 8'h8;
        my_rom[1280] = 8'h8;
        my_rom[1281] = 8'h8;
        my_rom[1282] = 8'h8;
        my_rom[1283] = 8'h8;
        my_rom[1284] = 8'h8;
        my_rom[1285] = 8'h8;
        my_rom[1286] = 8'h8;
        my_rom[1287] = 8'h8;
        my_rom[1288] = 8'ha;
        my_rom[1289] = 8'h8;
        my_rom[1290] = 8'h8;
        my_rom[1291] = 8'h8;
        my_rom[1292] = 8'h8;
        my_rom[1293] = 8'h8;
        my_rom[1294] = 8'h8;
        my_rom[1295] = 8'h8;
        my_rom[1296] = 8'h8;
        my_rom[1297] = 8'h8;
        my_rom[1298] = 8'h8;
        my_rom[1299] = 8'h8;
        my_rom[1300] = 8'h8;
        my_rom[1301] = 8'h8;
        my_rom[1302] = 8'h8;
        my_rom[1303] = 8'h8;
        my_rom[1304] = 8'h8;
        my_rom[1305] = 8'h8;
        my_rom[1306] = 8'h8;
        my_rom[1307] = 8'h8;
        my_rom[1308] = 8'h8;
        my_rom[1309] = 8'h8;
        my_rom[1310] = 8'h8;
        my_rom[1311] = 8'h8;
        my_rom[1312] = 8'h8;
        my_rom[1313] = 8'h8;
        my_rom[1314] = 8'h8;
        my_rom[1315] = 8'h8;
        my_rom[1316] = 8'h8;
        my_rom[1317] = 8'h8;
        my_rom[1318] = 8'h8;
        my_rom[1319] = 8'ha;
        my_rom[1320] = 8'h8;
        my_rom[1321] = 8'h8;
        my_rom[1322] = 8'h8;
        my_rom[1323] = 8'h8;
        my_rom[1324] = 8'h8;
        my_rom[1325] = 8'h8;
        my_rom[1326] = 8'h8;
        my_rom[1327] = 8'h8;
        my_rom[1328] = 8'h8;
        my_rom[1329] = 8'h8;
        my_rom[1330] = 8'h8;
        my_rom[1331] = 8'h8;
        my_rom[1332] = 8'h8;
        my_rom[1333] = 8'h8;
        my_rom[1334] = 8'h8;
        my_rom[1335] = 8'h8;
        my_rom[1336] = 8'h8;
        my_rom[1337] = 8'h8;
        my_rom[1338] = 8'h8;
        my_rom[1339] = 8'h8;
        my_rom[1340] = 8'h8;
        my_rom[1341] = 8'h8;
        my_rom[1342] = 8'h8;
        my_rom[1343] = 8'h8;
        my_rom[1344] = 8'h8;
        my_rom[1345] = 8'h8;
        my_rom[1346] = 8'h8;
        my_rom[1347] = 8'h8;
        my_rom[1348] = 8'h8;
        my_rom[1349] = 8'h8;
        my_rom[1350] = 8'ha;
        my_rom[1351] = 8'h8;
        my_rom[1352] = 8'h8;
        my_rom[1353] = 8'h8;
        my_rom[1354] = 8'h8;
        my_rom[1355] = 8'h8;
        my_rom[1356] = 8'h8;
        my_rom[1357] = 8'h8;
        my_rom[1358] = 8'h8;
        my_rom[1359] = 8'h8;
        my_rom[1360] = 8'h8;
        my_rom[1361] = 8'h8;
        my_rom[1362] = 8'h8;
        my_rom[1363] = 8'h8;
        my_rom[1364] = 8'h8;
        my_rom[1365] = 8'h8;
        my_rom[1366] = 8'h8;
        my_rom[1367] = 8'h8;
        my_rom[1368] = 8'h8;
        my_rom[1369] = 8'h8;
        my_rom[1370] = 8'h8;
        my_rom[1371] = 8'h8;
        my_rom[1372] = 8'h8;
        my_rom[1373] = 8'h8;
        my_rom[1374] = 8'h8;
        my_rom[1375] = 8'h8;
        my_rom[1376] = 8'h8;
        my_rom[1377] = 8'h8;
        my_rom[1378] = 8'h8;
        my_rom[1379] = 8'h8;
        my_rom[1380] = 8'h8;
        my_rom[1381] = 8'ha;
        my_rom[1382] = 8'h8;
        my_rom[1383] = 8'h8;
        my_rom[1384] = 8'h8;
        my_rom[1385] = 8'h8;
        my_rom[1386] = 8'h8;
        my_rom[1387] = 8'h8;
        my_rom[1388] = 8'h8;
        my_rom[1389] = 8'h8;
        my_rom[1390] = 8'h8;
        my_rom[1391] = 8'h8;
        my_rom[1392] = 8'h8;
        my_rom[1393] = 8'h8;
        my_rom[1394] = 8'h8;
        my_rom[1395] = 8'h8;
        my_rom[1396] = 8'h8;
        my_rom[1397] = 8'h8;
        my_rom[1398] = 8'h8;
        my_rom[1399] = 8'h8;
        my_rom[1400] = 8'h8;
        my_rom[1401] = 8'h8;
        my_rom[1402] = 8'h8;
        my_rom[1403] = 8'h8;
        my_rom[1404] = 8'h8;
        my_rom[1405] = 8'h8;
        my_rom[1406] = 8'h8;
        my_rom[1407] = 8'h8;
        my_rom[1408] = 8'h8;
        my_rom[1409] = 8'h8;
        my_rom[1410] = 8'h8;
        my_rom[1411] = 8'h8;
        my_rom[1412] = 8'ha;
        my_rom[1413] = 8'h8;
        my_rom[1414] = 8'h8;
        my_rom[1415] = 8'h8;
        my_rom[1416] = 8'h8;
        my_rom[1417] = 8'h8;
        my_rom[1418] = 8'h8;
        my_rom[1419] = 8'h8;
        my_rom[1420] = 8'h8;
        my_rom[1421] = 8'h8;
        my_rom[1422] = 8'h8;
        my_rom[1423] = 8'h8;
        my_rom[1424] = 8'h8;
        my_rom[1425] = 8'h8;
        my_rom[1426] = 8'h8;
        my_rom[1427] = 8'h8;
        my_rom[1428] = 8'h8;
        my_rom[1429] = 8'h8;
        my_rom[1430] = 8'h8;
        my_rom[1431] = 8'h8;
        my_rom[1432] = 8'h8;
        my_rom[1433] = 8'h8;
        my_rom[1434] = 8'h8;
        my_rom[1435] = 8'h8;
        my_rom[1436] = 8'h8;
        my_rom[1437] = 8'h8;
        my_rom[1438] = 8'h8;
        my_rom[1439] = 8'h8;
        my_rom[1440] = 8'h8;
        my_rom[1441] = 8'h8;
        my_rom[1442] = 8'h8;
        my_rom[1443] = 8'ha;
        my_rom[1444] = 8'h8;
        my_rom[1445] = 8'h8;
        my_rom[1446] = 8'h8;
        my_rom[1447] = 8'h8;
        my_rom[1448] = 8'h8;
        my_rom[1449] = 8'h8;
        my_rom[1450] = 8'h8;
        my_rom[1451] = 8'h8;
        my_rom[1452] = 8'h8;
        my_rom[1453] = 8'h8;
        my_rom[1454] = 8'h8;
        my_rom[1455] = 8'h8;
        my_rom[1456] = 8'h8;
        my_rom[1457] = 8'h8;
        my_rom[1458] = 8'h8;
        my_rom[1459] = 8'h8;
        my_rom[1460] = 8'h8;
        my_rom[1461] = 8'h8;
        my_rom[1462] = 8'h8;
        my_rom[1463] = 8'h8;
        my_rom[1464] = 8'h8;
        my_rom[1465] = 8'h8;
        my_rom[1466] = 8'h8;
        my_rom[1467] = 8'h8;
        my_rom[1468] = 8'h8;
        my_rom[1469] = 8'h8;
        my_rom[1470] = 8'h8;
        my_rom[1471] = 8'h8;
        my_rom[1472] = 8'h8;
        my_rom[1473] = 8'h8;
        my_rom[1474] = 8'ha;
        my_rom[1475] = 8'h8;
        my_rom[1476] = 8'h8;
        my_rom[1477] = 8'h8;
        my_rom[1478] = 8'h8;
        my_rom[1479] = 8'h8;
        my_rom[1480] = 8'h8;
        my_rom[1481] = 8'h8;
        my_rom[1482] = 8'h8;
        my_rom[1483] = 8'h8;
        my_rom[1484] = 8'h8;
        my_rom[1485] = 8'h8;
        my_rom[1486] = 8'h8;
        my_rom[1487] = 8'h8;
        my_rom[1488] = 8'h8;
        my_rom[1489] = 8'h8;
        my_rom[1490] = 8'h8;
        my_rom[1491] = 8'h8;
        my_rom[1492] = 8'h8;
        my_rom[1493] = 8'h8;
        my_rom[1494] = 8'h8;
        my_rom[1495] = 8'h8;
        my_rom[1496] = 8'h8;
        my_rom[1497] = 8'h8;
        my_rom[1498] = 8'h8;
        my_rom[1499] = 8'h8;
        my_rom[1500] = 8'h8;
        my_rom[1501] = 8'h8;
        my_rom[1502] = 8'h8;
        my_rom[1503] = 8'h8;
        my_rom[1504] = 8'h8;
        my_rom[1505] = 8'ha;
        my_rom[1506] = 8'h8;
        my_rom[1507] = 8'h8;
        my_rom[1508] = 8'h8;
        my_rom[1509] = 8'h8;
        my_rom[1510] = 8'h8;
        my_rom[1511] = 8'h8;
        my_rom[1512] = 8'h8;
        my_rom[1513] = 8'h8;
        my_rom[1514] = 8'h8;
        my_rom[1515] = 8'h8;
        my_rom[1516] = 8'h8;
        my_rom[1517] = 8'h8;
        my_rom[1518] = 8'h8;
        my_rom[1519] = 8'h8;
        my_rom[1520] = 8'h8;
        my_rom[1521] = 8'h8;
        my_rom[1522] = 8'h8;
        my_rom[1523] = 8'h8;
        my_rom[1524] = 8'h8;
        my_rom[1525] = 8'h8;
        my_rom[1526] = 8'h8;
        my_rom[1527] = 8'h8;
        my_rom[1528] = 8'h8;
        my_rom[1529] = 8'h8;
        my_rom[1530] = 8'h8;
        my_rom[1531] = 8'h8;
        my_rom[1532] = 8'h8;
        my_rom[1533] = 8'h8;
        my_rom[1534] = 8'h8;
        my_rom[1535] = 8'h8;
        my_rom[1536] = 8'ha;
        my_rom[1537] = 8'h8;
        my_rom[1538] = 8'h8;
        my_rom[1539] = 8'h8;
        my_rom[1540] = 8'h8;
        my_rom[1541] = 8'h8;
        my_rom[1542] = 8'h8;
        my_rom[1543] = 8'h8;
        my_rom[1544] = 8'h8;
        my_rom[1545] = 8'h8;
        my_rom[1546] = 8'h8;
        my_rom[1547] = 8'h8;
        my_rom[1548] = 8'h8;
        my_rom[1549] = 8'h8;
        my_rom[1550] = 8'h8;
        my_rom[1551] = 8'h8;
        my_rom[1552] = 8'h8;
        my_rom[1553] = 8'h8;
        my_rom[1554] = 8'h8;
        my_rom[1555] = 8'h8;
        my_rom[1556] = 8'h8;
        my_rom[1557] = 8'h8;
        my_rom[1558] = 8'h8;
        my_rom[1559] = 8'h8;
        my_rom[1560] = 8'h8;
        my_rom[1561] = 8'h8;
        my_rom[1562] = 8'h8;
        my_rom[1563] = 8'h8;
        my_rom[1564] = 8'h8;
        my_rom[1565] = 8'h8;
        my_rom[1566] = 8'h8;
        my_rom[1567] = 8'ha;
        my_rom[1568] = 8'h8;
        my_rom[1569] = 8'h8;
        my_rom[1570] = 8'h8;
        my_rom[1571] = 8'h8;
        my_rom[1572] = 8'h8;
        my_rom[1573] = 8'h8;
        my_rom[1574] = 8'h8;
        my_rom[1575] = 8'h8;
        my_rom[1576] = 8'h8;
        my_rom[1577] = 8'h8;
        my_rom[1578] = 8'h8;
        my_rom[1579] = 8'h8;
        my_rom[1580] = 8'h8;
        my_rom[1581] = 8'h8;
        my_rom[1582] = 8'h8;
        my_rom[1583] = 8'h8;
        my_rom[1584] = 8'h8;
        my_rom[1585] = 8'h8;
        my_rom[1586] = 8'h8;
        my_rom[1587] = 8'h8;
        my_rom[1588] = 8'h8;
        my_rom[1589] = 8'h8;
        my_rom[1590] = 8'h8;
        my_rom[1591] = 8'h8;
        my_rom[1592] = 8'h8;
        my_rom[1593] = 8'h8;
        my_rom[1594] = 8'h8;
        my_rom[1595] = 8'h8;
        my_rom[1596] = 8'h8;
        my_rom[1597] = 8'h8;
        my_rom[1598] = 8'ha;
        my_rom[1599] = 8'h8;
        my_rom[1600] = 8'h8;
        my_rom[1601] = 8'h8;
        my_rom[1602] = 8'h8;
        my_rom[1603] = 8'h8;
        my_rom[1604] = 8'h8;
        my_rom[1605] = 8'h8;
        my_rom[1606] = 8'h8;
        my_rom[1607] = 8'h8;
        my_rom[1608] = 8'h8;
        my_rom[1609] = 8'h8;
        my_rom[1610] = 8'h8;
        my_rom[1611] = 8'h8;
        my_rom[1612] = 8'h8;
        my_rom[1613] = 8'h8;
        my_rom[1614] = 8'h8;
        my_rom[1615] = 8'h8;
        my_rom[1616] = 8'h8;
        my_rom[1617] = 8'h8;
        my_rom[1618] = 8'h8;
        my_rom[1619] = 8'h8;
        my_rom[1620] = 8'h8;
        my_rom[1621] = 8'h8;
        my_rom[1622] = 8'h8;
        my_rom[1623] = 8'h8;
        my_rom[1624] = 8'h8;
        my_rom[1625] = 8'h8;
        my_rom[1626] = 8'h8;
        my_rom[1627] = 8'h8;
        my_rom[1628] = 8'h8;
        my_rom[1629] = 8'ha;
        my_rom[1630] = 8'hc;
        my_rom[1631] = 8'h0;
        my_rom[1632] = 8'h8;
        my_rom[1633] = 8'h8;
        my_rom[1634] = 8'h8;
        my_rom[1635] = 8'h8;
        my_rom[1636] = 8'h8;
        my_rom[1637] = 8'h8;
        my_rom[1638] = 8'h8;
        my_rom[1639] = 8'h8;
        my_rom[1640] = 8'h8;
        my_rom[1641] = 8'h8;
        my_rom[1642] = 8'h8;
        my_rom[1643] = 8'h8;
        my_rom[1644] = 8'h8;
        my_rom[1645] = 8'h8;
        my_rom[1646] = 8'h8;
        my_rom[1647] = 8'h8;
        my_rom[1648] = 8'h8;
        my_rom[1649] = 8'h8;
        my_rom[1650] = 8'h8;
        my_rom[1651] = 8'h8;
        my_rom[1652] = 8'h8;
        my_rom[1653] = 8'h8;
        my_rom[1654] = 8'h8;
        my_rom[1655] = 8'h8;
        my_rom[1656] = 8'h8;
        my_rom[1657] = 8'h8;
        my_rom[1658] = 8'h8;
        my_rom[1659] = 8'h8;
        my_rom[1660] = 8'h8;
        my_rom[1661] = 8'h8;
        my_rom[1662] = 8'hf5;
        my_rom[1663] = 8'hf5;
        my_rom[1664] = 8'ha5;
        my_rom[1665] = 8'ha5;
        my_rom[1666] = 8'ha5;
        my_rom[1667] = 8'ha5;
        my_rom[1668] = 8'had;
        my_rom[1669] = 8'had;
        my_rom[1670] = 8'ha5;
        my_rom[1671] = 8'had;
        my_rom[1672] = 8'had;
        my_rom[1673] = 8'h8;
        my_rom[1674] = 8'h8;
        my_rom[1675] = 8'h8;
        my_rom[1676] = 8'h8;
        my_rom[1677] = 8'h8;
        my_rom[1678] = 8'h8;
        my_rom[1679] = 8'h8;
        my_rom[1680] = 8'h8;
        my_rom[1681] = 8'h8;
        my_rom[1682] = 8'h8;
        my_rom[1683] = 8'h8;
        my_rom[1684] = 8'h8;
        my_rom[1685] = 8'h8;
        my_rom[1686] = 8'h8;
        my_rom[1687] = 8'h8;
        my_rom[1688] = 8'h8;
        my_rom[1689] = 8'h8;
        my_rom[1690] = 8'h8;
        my_rom[1691] = 8'ha;
        my_rom[1692] = 8'h8;
        my_rom[1693] = 8'h8;
        my_rom[1694] = 8'h8;
        my_rom[1695] = 8'h8;
        my_rom[1696] = 8'h8;
        my_rom[1697] = 8'h8;
        my_rom[1698] = 8'h8;
        my_rom[1699] = 8'h8;
        my_rom[1700] = 8'h8;
        my_rom[1701] = 8'h8;
        my_rom[1702] = 8'h8;
        my_rom[1703] = 8'h8;
        my_rom[1704] = 8'h8;
        my_rom[1705] = 8'h8;
        my_rom[1706] = 8'h8;
        my_rom[1707] = 8'h8;
        my_rom[1708] = 8'h8;
        my_rom[1709] = 8'h8;
        my_rom[1710] = 8'h8;
        my_rom[1711] = 8'h8;
        my_rom[1712] = 8'h8;
        my_rom[1713] = 8'h8;
        my_rom[1714] = 8'hf5;
        my_rom[1715] = 8'had;
        my_rom[1716] = 8'had;
        my_rom[1717] = 8'hed;
        my_rom[1718] = 8'hed;
        my_rom[1719] = 8'had;
        my_rom[1720] = 8'ha5;
        my_rom[1721] = 8'ha5;
        my_rom[1722] = 8'ha5;
        my_rom[1723] = 8'ha5;
        my_rom[1724] = 8'ha5;
        my_rom[1725] = 8'h9d;
        my_rom[1726] = 8'h9b;
        my_rom[1727] = 8'ha5;
        my_rom[1728] = 8'ha5;
        my_rom[1729] = 8'ha5;
        my_rom[1730] = 8'ha5;
        my_rom[1731] = 8'ha5;
        my_rom[1732] = 8'ha5;
        my_rom[1733] = 8'ha5;
        my_rom[1734] = 8'h5b;
        my_rom[1735] = 8'h53;
        my_rom[1736] = 8'h8;
        my_rom[1737] = 8'h8;
        my_rom[1738] = 8'h8;
        my_rom[1739] = 8'h8;
        my_rom[1740] = 8'h8;
        my_rom[1741] = 8'h8;
        my_rom[1742] = 8'h8;
        my_rom[1743] = 8'h8;
        my_rom[1744] = 8'h8;
        my_rom[1745] = 8'h8;
        my_rom[1746] = 8'h8;
        my_rom[1747] = 8'h8;
        my_rom[1748] = 8'h8;
        my_rom[1749] = 8'h8;
        my_rom[1750] = 8'h8;
        my_rom[1751] = 8'ha;
        my_rom[1752] = 8'h8;
        my_rom[1753] = 8'h8;
        my_rom[1754] = 8'h8;
        my_rom[1755] = 8'h8;
        my_rom[1756] = 8'h8;
        my_rom[1757] = 8'h8;
        my_rom[1758] = 8'h8;
        my_rom[1759] = 8'h8;
        my_rom[1760] = 8'h8;
        my_rom[1761] = 8'h8;
        my_rom[1762] = 8'h8;
        my_rom[1763] = 8'h8;
        my_rom[1764] = 8'h8;
        my_rom[1765] = 8'h8;
        my_rom[1766] = 8'h8;
        my_rom[1767] = 8'h8;
        my_rom[1768] = 8'h8;
        my_rom[1769] = 8'h8;
        my_rom[1770] = 8'had;
        my_rom[1771] = 8'had;
        my_rom[1772] = 8'hf5;
        my_rom[1773] = 8'hf5;
        my_rom[1774] = 8'hed;
        my_rom[1775] = 8'ha5;
        my_rom[1776] = 8'ha5;
        my_rom[1777] = 8'ha5;
        my_rom[1778] = 8'ha5;
        my_rom[1779] = 8'h9d;
        my_rom[1780] = 8'h9b;
        my_rom[1781] = 8'h5b;
        my_rom[1782] = 8'h9b;
        my_rom[1783] = 8'h5b;
        my_rom[1784] = 8'h5b;
        my_rom[1785] = 8'h5b;
        my_rom[1786] = 8'h9b;
        my_rom[1787] = 8'h9d;
        my_rom[1788] = 8'h9d;
        my_rom[1789] = 8'ha5;
        my_rom[1790] = 8'ha5;
        my_rom[1791] = 8'ha5;
        my_rom[1792] = 8'ha5;
        my_rom[1793] = 8'ha5;
        my_rom[1794] = 8'h5b;
        my_rom[1795] = 8'h53;
        my_rom[1796] = 8'h8;
        my_rom[1797] = 8'h8;
        my_rom[1798] = 8'h8;
        my_rom[1799] = 8'h8;
        my_rom[1800] = 8'h8;
        my_rom[1801] = 8'h8;
        my_rom[1802] = 8'h8;
        my_rom[1803] = 8'h8;
        my_rom[1804] = 8'h8;
        my_rom[1805] = 8'h8;
        my_rom[1806] = 8'h8;
        my_rom[1807] = 8'h8;
        my_rom[1808] = 8'h8;
        my_rom[1809] = 8'h8;
        my_rom[1810] = 8'h8;
        my_rom[1811] = 8'ha;
        my_rom[1812] = 8'h8;
        my_rom[1813] = 8'h8;
        my_rom[1814] = 8'h8;
        my_rom[1815] = 8'h8;
        my_rom[1816] = 8'h8;
        my_rom[1817] = 8'h8;
        my_rom[1818] = 8'h8;
        my_rom[1819] = 8'h8;
        my_rom[1820] = 8'h8;
        my_rom[1821] = 8'h8;
        my_rom[1822] = 8'h8;
        my_rom[1823] = 8'h8;
        my_rom[1824] = 8'h8;
        my_rom[1825] = 8'h8;
        my_rom[1826] = 8'h8;
        my_rom[1827] = 8'ha3;
        my_rom[1828] = 8'ha5;
        my_rom[1829] = 8'ha5;
        my_rom[1830] = 8'ha5;
        my_rom[1831] = 8'had;
        my_rom[1832] = 8'ha5;
        my_rom[1833] = 8'ha5;
        my_rom[1834] = 8'ha5;
        my_rom[1835] = 8'ha5;
        my_rom[1836] = 8'h9d;
        my_rom[1837] = 8'ha5;
        my_rom[1838] = 8'h9d;
        my_rom[1839] = 8'h5b;
        my_rom[1840] = 8'h5b;
        my_rom[1841] = 8'h5b;
        my_rom[1842] = 8'h5b;
        my_rom[1843] = 8'h5b;
        my_rom[1844] = 8'h5b;
        my_rom[1845] = 8'h53;
        my_rom[1846] = 8'h53;
        my_rom[1847] = 8'h53;
        my_rom[1848] = 8'h53;
        my_rom[1849] = 8'h53;
        my_rom[1850] = 8'h5b;
        my_rom[1851] = 8'h9d;
        my_rom[1852] = 8'ha5;
        my_rom[1853] = 8'ha5;
        my_rom[1854] = 8'h5b;
        my_rom[1855] = 8'h5b;
        my_rom[1856] = 8'h53;
        my_rom[1857] = 8'h8;
        my_rom[1858] = 8'h8;
        my_rom[1859] = 8'h8;
        my_rom[1860] = 8'h8;
        my_rom[1861] = 8'h8;
        my_rom[1862] = 8'h8;
        my_rom[1863] = 8'h8;
        my_rom[1864] = 8'h8;
        my_rom[1865] = 8'h8;
        my_rom[1866] = 8'h8;
        my_rom[1867] = 8'h8;
        my_rom[1868] = 8'h8;
        my_rom[1869] = 8'h8;
        my_rom[1870] = 8'h8;
        my_rom[1871] = 8'ha;
        my_rom[1872] = 8'h8;
        my_rom[1873] = 8'h8;
        my_rom[1874] = 8'h8;
        my_rom[1875] = 8'h8;
        my_rom[1876] = 8'h8;
        my_rom[1877] = 8'h8;
        my_rom[1878] = 8'h8;
        my_rom[1879] = 8'h8;
        my_rom[1880] = 8'h8;
        my_rom[1881] = 8'h8;
        my_rom[1882] = 8'h8;
        my_rom[1883] = 8'h8;
        my_rom[1884] = 8'h8;
        my_rom[1885] = 8'h8;
        my_rom[1886] = 8'ha3;
        my_rom[1887] = 8'ha5;
        my_rom[1888] = 8'ha3;
        my_rom[1889] = 8'h9b;
        my_rom[1890] = 8'h9b;
        my_rom[1891] = 8'h9b;
        my_rom[1892] = 8'h9b;
        my_rom[1893] = 8'ha5;
        my_rom[1894] = 8'ha5;
        my_rom[1895] = 8'h9d;
        my_rom[1896] = 8'h9b;
        my_rom[1897] = 8'h9d;
        my_rom[1898] = 8'h5b;
        my_rom[1899] = 8'h5b;
        my_rom[1900] = 8'h5b;
        my_rom[1901] = 8'h5b;
        my_rom[1902] = 8'h53;
        my_rom[1903] = 8'h53;
        my_rom[1904] = 8'h53;
        my_rom[1905] = 8'h53;
        my_rom[1906] = 8'h53;
        my_rom[1907] = 8'h4b;
        my_rom[1908] = 8'h4b;
        my_rom[1909] = 8'h53;
        my_rom[1910] = 8'h53;
        my_rom[1911] = 8'h53;
        my_rom[1912] = 8'h53;
        my_rom[1913] = 8'h5b;
        my_rom[1914] = 8'h9b;
        my_rom[1915] = 8'h5b;
        my_rom[1916] = 8'h5b;
        my_rom[1917] = 8'h8;
        my_rom[1918] = 8'h8;
        my_rom[1919] = 8'h8;
        my_rom[1920] = 8'h8;
        my_rom[1921] = 8'h8;
        my_rom[1922] = 8'h8;
        my_rom[1923] = 8'h8;
        my_rom[1924] = 8'h8;
        my_rom[1925] = 8'h8;
        my_rom[1926] = 8'h8;
        my_rom[1927] = 8'h8;
        my_rom[1928] = 8'h8;
        my_rom[1929] = 8'h8;
        my_rom[1930] = 8'h8;
        my_rom[1931] = 8'ha;
        my_rom[1932] = 8'h8;
        my_rom[1933] = 8'h8;
        my_rom[1934] = 8'h8;
        my_rom[1935] = 8'h8;
        my_rom[1936] = 8'h8;
        my_rom[1937] = 8'h8;
        my_rom[1938] = 8'h8;
        my_rom[1939] = 8'h8;
        my_rom[1940] = 8'h8;
        my_rom[1941] = 8'h8;
        my_rom[1942] = 8'h8;
        my_rom[1943] = 8'h8;
        my_rom[1944] = 8'h8;
        my_rom[1945] = 8'ha3;
        my_rom[1946] = 8'ha3;
        my_rom[1947] = 8'h9b;
        my_rom[1948] = 8'h9b;
        my_rom[1949] = 8'h5b;
        my_rom[1950] = 8'h5b;
        my_rom[1951] = 8'h9b;
        my_rom[1952] = 8'h9b;
        my_rom[1953] = 8'ha3;
        my_rom[1954] = 8'h9b;
        my_rom[1955] = 8'h9b;
        my_rom[1956] = 8'h9b;
        my_rom[1957] = 8'h9b;
        my_rom[1958] = 8'h9b;
        my_rom[1959] = 8'h5b;
        my_rom[1960] = 8'h5b;
        my_rom[1961] = 8'h53;
        my_rom[1962] = 8'h53;
        my_rom[1963] = 8'hb;
        my_rom[1964] = 8'hb;
        my_rom[1965] = 8'hb;
        my_rom[1966] = 8'h53;
        my_rom[1967] = 8'h53;
        my_rom[1968] = 8'h53;
        my_rom[1969] = 8'h53;
        my_rom[1970] = 8'h53;
        my_rom[1971] = 8'h53;
        my_rom[1972] = 8'h53;
        my_rom[1973] = 8'h53;
        my_rom[1974] = 8'h5b;
        my_rom[1975] = 8'h5b;
        my_rom[1976] = 8'h53;
        my_rom[1977] = 8'h53;
        my_rom[1978] = 8'h53;
        my_rom[1979] = 8'h8;
        my_rom[1980] = 8'h8;
        my_rom[1981] = 8'h8;
        my_rom[1982] = 8'h8;
        my_rom[1983] = 8'h8;
        my_rom[1984] = 8'h8;
        my_rom[1985] = 8'h8;
        my_rom[1986] = 8'h8;
        my_rom[1987] = 8'h8;
        my_rom[1988] = 8'h8;
        my_rom[1989] = 8'h8;
        my_rom[1990] = 8'h8;
        my_rom[1991] = 8'ha;
        my_rom[1992] = 8'h8;
        my_rom[1993] = 8'h8;
        my_rom[1994] = 8'h8;
        my_rom[1995] = 8'h8;
        my_rom[1996] = 8'h8;
        my_rom[1997] = 8'h8;
        my_rom[1998] = 8'h8;
        my_rom[1999] = 8'h8;
        my_rom[2000] = 8'h8;
        my_rom[2001] = 8'h8;
        my_rom[2002] = 8'h8;
        my_rom[2003] = 8'h8;
        my_rom[2004] = 8'h9b;
        my_rom[2005] = 8'h9b;
        my_rom[2006] = 8'h9b;
        my_rom[2007] = 8'h5b;
        my_rom[2008] = 8'h5b;
        my_rom[2009] = 8'h53;
        my_rom[2010] = 8'h5b;
        my_rom[2011] = 8'h9b;
        my_rom[2012] = 8'h9b;
        my_rom[2013] = 8'h9b;
        my_rom[2014] = 8'h9b;
        my_rom[2015] = 8'h9b;
        my_rom[2016] = 8'h9b;
        my_rom[2017] = 8'h5b;
        my_rom[2018] = 8'h53;
        my_rom[2019] = 8'h5b;
        my_rom[2020] = 8'h5b;
        my_rom[2021] = 8'h53;
        my_rom[2022] = 8'h53;
        my_rom[2023] = 8'h53;
        my_rom[2024] = 8'h53;
        my_rom[2025] = 8'h53;
        my_rom[2026] = 8'h53;
        my_rom[2027] = 8'h53;
        my_rom[2028] = 8'h53;
        my_rom[2029] = 8'h53;
        my_rom[2030] = 8'h53;
        my_rom[2031] = 8'h53;
        my_rom[2032] = 8'h53;
        my_rom[2033] = 8'h53;
        my_rom[2034] = 8'h53;
        my_rom[2035] = 8'h53;
        my_rom[2036] = 8'h5b;
        my_rom[2037] = 8'h5b;
        my_rom[2038] = 8'h5b;
        my_rom[2039] = 8'h5b;
        my_rom[2040] = 8'h8;
        my_rom[2041] = 8'h8;
        my_rom[2042] = 8'h8;
        my_rom[2043] = 8'h8;
        my_rom[2044] = 8'h8;
        my_rom[2045] = 8'h8;
        my_rom[2046] = 8'h8;
        my_rom[2047] = 8'h8;
        my_rom[2048] = 8'h8;
        my_rom[2049] = 8'h8;
        my_rom[2050] = 8'h8;
        my_rom[2051] = 8'ha;
        my_rom[2052] = 8'h8;
        my_rom[2053] = 8'h8;
        my_rom[2054] = 8'h8;
        my_rom[2055] = 8'h8;
        my_rom[2056] = 8'h8;
        my_rom[2057] = 8'h8;
        my_rom[2058] = 8'h8;
        my_rom[2059] = 8'h8;
        my_rom[2060] = 8'h8;
        my_rom[2061] = 8'h8;
        my_rom[2062] = 8'h8;
        my_rom[2063] = 8'ha3;
        my_rom[2064] = 8'ha3;
        my_rom[2065] = 8'h9b;
        my_rom[2066] = 8'h5b;
        my_rom[2067] = 8'h53;
        my_rom[2068] = 8'h53;
        my_rom[2069] = 8'h53;
        my_rom[2070] = 8'h53;
        my_rom[2071] = 8'h9b;
        my_rom[2072] = 8'h53;
        my_rom[2073] = 8'h53;
        my_rom[2074] = 8'h53;
        my_rom[2075] = 8'h53;
        my_rom[2076] = 8'h5b;
        my_rom[2077] = 8'h9b;
        my_rom[2078] = 8'h9b;
        my_rom[2079] = 8'h53;
        my_rom[2080] = 8'h53;
        my_rom[2081] = 8'h53;
        my_rom[2082] = 8'h53;
        my_rom[2083] = 8'h53;
        my_rom[2084] = 8'h53;
        my_rom[2085] = 8'h53;
        my_rom[2086] = 8'h53;
        my_rom[2087] = 8'h53;
        my_rom[2088] = 8'h53;
        my_rom[2089] = 8'h53;
        my_rom[2090] = 8'h53;
        my_rom[2091] = 8'h53;
        my_rom[2092] = 8'h53;
        my_rom[2093] = 8'h53;
        my_rom[2094] = 8'h53;
        my_rom[2095] = 8'h53;
        my_rom[2096] = 8'h53;
        my_rom[2097] = 8'h5b;
        my_rom[2098] = 8'h5b;
        my_rom[2099] = 8'h5b;
        my_rom[2100] = 8'h5b;
        my_rom[2101] = 8'h8;
        my_rom[2102] = 8'h8;
        my_rom[2103] = 8'h8;
        my_rom[2104] = 8'h8;
        my_rom[2105] = 8'h8;
        my_rom[2106] = 8'h8;
        my_rom[2107] = 8'h8;
        my_rom[2108] = 8'h8;
        my_rom[2109] = 8'h8;
        my_rom[2110] = 8'h8;
        my_rom[2111] = 8'ha;
        my_rom[2112] = 8'h8;
        my_rom[2113] = 8'h8;
        my_rom[2114] = 8'h8;
        my_rom[2115] = 8'h8;
        my_rom[2116] = 8'h8;
        my_rom[2117] = 8'h8;
        my_rom[2118] = 8'h8;
        my_rom[2119] = 8'h8;
        my_rom[2120] = 8'h8;
        my_rom[2121] = 8'h8;
        my_rom[2122] = 8'ha5;
        my_rom[2123] = 8'ha3;
        my_rom[2124] = 8'h5b;
        my_rom[2125] = 8'h5b;
        my_rom[2126] = 8'h53;
        my_rom[2127] = 8'h53;
        my_rom[2128] = 8'h53;
        my_rom[2129] = 8'h53;
        my_rom[2130] = 8'h53;
        my_rom[2131] = 8'h53;
        my_rom[2132] = 8'h53;
        my_rom[2133] = 8'h49;
        my_rom[2134] = 8'h4b;
        my_rom[2135] = 8'h53;
        my_rom[2136] = 8'h53;
        my_rom[2137] = 8'h53;
        my_rom[2138] = 8'h53;
        my_rom[2139] = 8'h53;
        my_rom[2140] = 8'h53;
        my_rom[2141] = 8'h53;
        my_rom[2142] = 8'h53;
        my_rom[2143] = 8'h53;
        my_rom[2144] = 8'h53;
        my_rom[2145] = 8'h53;
        my_rom[2146] = 8'h53;
        my_rom[2147] = 8'h53;
        my_rom[2148] = 8'h4b;
        my_rom[2149] = 8'hb;
        my_rom[2150] = 8'hb;
        my_rom[2151] = 8'hb;
        my_rom[2152] = 8'hb;
        my_rom[2153] = 8'h4b;
        my_rom[2154] = 8'h4b;
        my_rom[2155] = 8'h53;
        my_rom[2156] = 8'h53;
        my_rom[2157] = 8'h53;
        my_rom[2158] = 8'h53;
        my_rom[2159] = 8'h5b;
        my_rom[2160] = 8'h5b;
        my_rom[2161] = 8'h8;
        my_rom[2162] = 8'h8;
        my_rom[2163] = 8'h8;
        my_rom[2164] = 8'h8;
        my_rom[2165] = 8'h8;
        my_rom[2166] = 8'h8;
        my_rom[2167] = 8'h8;
        my_rom[2168] = 8'h8;
        my_rom[2169] = 8'h8;
        my_rom[2170] = 8'h8;
        my_rom[2171] = 8'ha;
        my_rom[2172] = 8'h8;
        my_rom[2173] = 8'h8;
        my_rom[2174] = 8'h8;
        my_rom[2175] = 8'h8;
        my_rom[2176] = 8'h8;
        my_rom[2177] = 8'h8;
        my_rom[2178] = 8'h8;
        my_rom[2179] = 8'h8;
        my_rom[2180] = 8'h8;
        my_rom[2181] = 8'h8;
        my_rom[2182] = 8'ha5;
        my_rom[2183] = 8'h9b;
        my_rom[2184] = 8'h53;
        my_rom[2185] = 8'h53;
        my_rom[2186] = 8'h53;
        my_rom[2187] = 8'h53;
        my_rom[2188] = 8'h53;
        my_rom[2189] = 8'h53;
        my_rom[2190] = 8'h49;
        my_rom[2191] = 8'h9;
        my_rom[2192] = 8'h9;
        my_rom[2193] = 8'h9;
        my_rom[2194] = 8'h9;
        my_rom[2195] = 8'h9;
        my_rom[2196] = 8'h49;
        my_rom[2197] = 8'h49;
        my_rom[2198] = 8'h49;
        my_rom[2199] = 8'h53;
        my_rom[2200] = 8'h53;
        my_rom[2201] = 8'h53;
        my_rom[2202] = 8'h53;
        my_rom[2203] = 8'h53;
        my_rom[2204] = 8'h53;
        my_rom[2205] = 8'h53;
        my_rom[2206] = 8'h53;
        my_rom[2207] = 8'h4b;
        my_rom[2208] = 8'h53;
        my_rom[2209] = 8'hb;
        my_rom[2210] = 8'hb;
        my_rom[2211] = 8'hb;
        my_rom[2212] = 8'hb;
        my_rom[2213] = 8'hb;
        my_rom[2214] = 8'hb;
        my_rom[2215] = 8'hb;
        my_rom[2216] = 8'h4b;
        my_rom[2217] = 8'h53;
        my_rom[2218] = 8'h53;
        my_rom[2219] = 8'h53;
        my_rom[2220] = 8'h5b;
        my_rom[2221] = 8'h5b;
        my_rom[2222] = 8'h8;
        my_rom[2223] = 8'h8;
        my_rom[2224] = 8'h8;
        my_rom[2225] = 8'h8;
        my_rom[2226] = 8'h8;
        my_rom[2227] = 8'h8;
        my_rom[2228] = 8'h8;
        my_rom[2229] = 8'h8;
        my_rom[2230] = 8'h8;
        my_rom[2231] = 8'ha;
        my_rom[2232] = 8'h8;
        my_rom[2233] = 8'h8;
        my_rom[2234] = 8'h8;
        my_rom[2235] = 8'h8;
        my_rom[2236] = 8'h8;
        my_rom[2237] = 8'h8;
        my_rom[2238] = 8'h8;
        my_rom[2239] = 8'h8;
        my_rom[2240] = 8'ha5;
        my_rom[2241] = 8'ha5;
        my_rom[2242] = 8'h9b;
        my_rom[2243] = 8'h53;
        my_rom[2244] = 8'h53;
        my_rom[2245] = 8'h53;
        my_rom[2246] = 8'h53;
        my_rom[2247] = 8'h53;
        my_rom[2248] = 8'h49;
        my_rom[2249] = 8'h49;
        my_rom[2250] = 8'h9;
        my_rom[2251] = 8'h1;
        my_rom[2252] = 8'h1;
        my_rom[2253] = 8'h1;
        my_rom[2254] = 8'h9;
        my_rom[2255] = 8'h1;
        my_rom[2256] = 8'h1;
        my_rom[2257] = 8'h9;
        my_rom[2258] = 8'h53;
        my_rom[2259] = 8'h53;
        my_rom[2260] = 8'h53;
        my_rom[2261] = 8'h53;
        my_rom[2262] = 8'h53;
        my_rom[2263] = 8'h53;
        my_rom[2264] = 8'h53;
        my_rom[2265] = 8'h53;
        my_rom[2266] = 8'h4b;
        my_rom[2267] = 8'h4b;
        my_rom[2268] = 8'hb;
        my_rom[2269] = 8'hb;
        my_rom[2270] = 8'hb;
        my_rom[2271] = 8'hb;
        my_rom[2272] = 8'hb;
        my_rom[2273] = 8'hb;
        my_rom[2274] = 8'hb;
        my_rom[2275] = 8'hb;
        my_rom[2276] = 8'hb;
        my_rom[2277] = 8'hb;
        my_rom[2278] = 8'h53;
        my_rom[2279] = 8'h5b;
        my_rom[2280] = 8'h5b;
        my_rom[2281] = 8'h53;
        my_rom[2282] = 8'h53;
        my_rom[2283] = 8'h8;
        my_rom[2284] = 8'h8;
        my_rom[2285] = 8'h8;
        my_rom[2286] = 8'h8;
        my_rom[2287] = 8'h8;
        my_rom[2288] = 8'h8;
        my_rom[2289] = 8'h8;
        my_rom[2290] = 8'h8;
        my_rom[2291] = 8'ha;
        my_rom[2292] = 8'h8;
        my_rom[2293] = 8'h8;
        my_rom[2294] = 8'h8;
        my_rom[2295] = 8'h8;
        my_rom[2296] = 8'h8;
        my_rom[2297] = 8'h8;
        my_rom[2298] = 8'h8;
        my_rom[2299] = 8'h8;
        my_rom[2300] = 8'had;
        my_rom[2301] = 8'h9b;
        my_rom[2302] = 8'h5b;
        my_rom[2303] = 8'h53;
        my_rom[2304] = 8'h53;
        my_rom[2305] = 8'h53;
        my_rom[2306] = 8'h53;
        my_rom[2307] = 8'h49;
        my_rom[2308] = 8'h9;
        my_rom[2309] = 8'h49;
        my_rom[2310] = 8'h9;
        my_rom[2311] = 8'h9;
        my_rom[2312] = 8'h1;
        my_rom[2313] = 8'h1;
        my_rom[2314] = 8'h9;
        my_rom[2315] = 8'h1;
        my_rom[2316] = 8'h1;
        my_rom[2317] = 8'h9;
        my_rom[2318] = 8'h49;
        my_rom[2319] = 8'h53;
        my_rom[2320] = 8'h53;
        my_rom[2321] = 8'h53;
        my_rom[2322] = 8'h53;
        my_rom[2323] = 8'h53;
        my_rom[2324] = 8'h53;
        my_rom[2325] = 8'h4b;
        my_rom[2326] = 8'h9;
        my_rom[2327] = 8'h9;
        my_rom[2328] = 8'h9;
        my_rom[2329] = 8'h9;
        my_rom[2330] = 8'h9;
        my_rom[2331] = 8'hb;
        my_rom[2332] = 8'hb;
        my_rom[2333] = 8'hb;
        my_rom[2334] = 8'hb;
        my_rom[2335] = 8'hb;
        my_rom[2336] = 8'hb;
        my_rom[2337] = 8'h53;
        my_rom[2338] = 8'h4b;
        my_rom[2339] = 8'h53;
        my_rom[2340] = 8'h5b;
        my_rom[2341] = 8'h5b;
        my_rom[2342] = 8'h5b;
        my_rom[2343] = 8'h8;
        my_rom[2344] = 8'h8;
        my_rom[2345] = 8'h8;
        my_rom[2346] = 8'h8;
        my_rom[2347] = 8'h8;
        my_rom[2348] = 8'h8;
        my_rom[2349] = 8'h8;
        my_rom[2350] = 8'h8;
        my_rom[2351] = 8'ha;
        my_rom[2352] = 8'h8;
        my_rom[2353] = 8'h8;
        my_rom[2354] = 8'h8;
        my_rom[2355] = 8'h8;
        my_rom[2356] = 8'h8;
        my_rom[2357] = 8'h8;
        my_rom[2358] = 8'h8;
        my_rom[2359] = 8'had;
        my_rom[2360] = 8'ha5;
        my_rom[2361] = 8'h53;
        my_rom[2362] = 8'h53;
        my_rom[2363] = 8'h53;
        my_rom[2364] = 8'h53;
        my_rom[2365] = 8'h53;
        my_rom[2366] = 8'h53;
        my_rom[2367] = 8'h53;
        my_rom[2368] = 8'h49;
        my_rom[2369] = 8'h49;
        my_rom[2370] = 8'h49;
        my_rom[2371] = 8'h9;
        my_rom[2372] = 8'h9;
        my_rom[2373] = 8'h9;
        my_rom[2374] = 8'h49;
        my_rom[2375] = 8'h9;
        my_rom[2376] = 8'h9;
        my_rom[2377] = 8'h9;
        my_rom[2378] = 8'h1;
        my_rom[2379] = 8'h49;
        my_rom[2380] = 8'h5b;
        my_rom[2381] = 8'h9d;
        my_rom[2382] = 8'h5b;
        my_rom[2383] = 8'h53;
        my_rom[2384] = 8'h53;
        my_rom[2385] = 8'h4b;
        my_rom[2386] = 8'h4b;
        my_rom[2387] = 8'hb;
        my_rom[2388] = 8'hb;
        my_rom[2389] = 8'h9;
        my_rom[2390] = 8'h9;
        my_rom[2391] = 8'h9;
        my_rom[2392] = 8'h9;
        my_rom[2393] = 8'hb;
        my_rom[2394] = 8'hb;
        my_rom[2395] = 8'hb;
        my_rom[2396] = 8'hb;
        my_rom[2397] = 8'hb;
        my_rom[2398] = 8'h53;
        my_rom[2399] = 8'h53;
        my_rom[2400] = 8'h53;
        my_rom[2401] = 8'h5b;
        my_rom[2402] = 8'h5b;
        my_rom[2403] = 8'h8;
        my_rom[2404] = 8'h8;
        my_rom[2405] = 8'h8;
        my_rom[2406] = 8'h8;
        my_rom[2407] = 8'h8;
        my_rom[2408] = 8'h8;
        my_rom[2409] = 8'h8;
        my_rom[2410] = 8'h8;
        my_rom[2411] = 8'ha;
        my_rom[2412] = 8'h8;
        my_rom[2413] = 8'h8;
        my_rom[2414] = 8'h8;
        my_rom[2415] = 8'h8;
        my_rom[2416] = 8'h8;
        my_rom[2417] = 8'h8;
        my_rom[2418] = 8'h8;
        my_rom[2419] = 8'ha5;
        my_rom[2420] = 8'h53;
        my_rom[2421] = 8'h53;
        my_rom[2422] = 8'h53;
        my_rom[2423] = 8'h53;
        my_rom[2424] = 8'h53;
        my_rom[2425] = 8'h53;
        my_rom[2426] = 8'h53;
        my_rom[2427] = 8'h53;
        my_rom[2428] = 8'h53;
        my_rom[2429] = 8'h53;
        my_rom[2430] = 8'h53;
        my_rom[2431] = 8'h53;
        my_rom[2432] = 8'h53;
        my_rom[2433] = 8'h53;
        my_rom[2434] = 8'h53;
        my_rom[2435] = 8'h53;
        my_rom[2436] = 8'h53;
        my_rom[2437] = 8'h49;
        my_rom[2438] = 8'h49;
        my_rom[2439] = 8'h49;
        my_rom[2440] = 8'h49;
        my_rom[2441] = 8'h53;
        my_rom[2442] = 8'h53;
        my_rom[2443] = 8'h53;
        my_rom[2444] = 8'h4b;
        my_rom[2445] = 8'h4b;
        my_rom[2446] = 8'h9;
        my_rom[2447] = 8'h9;
        my_rom[2448] = 8'h9;
        my_rom[2449] = 8'h9;
        my_rom[2450] = 8'h9;
        my_rom[2451] = 8'h9;
        my_rom[2452] = 8'h9;
        my_rom[2453] = 8'h9;
        my_rom[2454] = 8'h9;
        my_rom[2455] = 8'h9;
        my_rom[2456] = 8'hb;
        my_rom[2457] = 8'hb;
        my_rom[2458] = 8'hb;
        my_rom[2459] = 8'h4b;
        my_rom[2460] = 8'h53;
        my_rom[2461] = 8'h53;
        my_rom[2462] = 8'h5b;
        my_rom[2463] = 8'h53;
        my_rom[2464] = 8'h8;
        my_rom[2465] = 8'h8;
        my_rom[2466] = 8'h8;
        my_rom[2467] = 8'h8;
        my_rom[2468] = 8'h8;
        my_rom[2469] = 8'h8;
        my_rom[2470] = 8'h8;
        my_rom[2471] = 8'ha;
        my_rom[2472] = 8'h8;
        my_rom[2473] = 8'h8;
        my_rom[2474] = 8'h8;
        my_rom[2475] = 8'h8;
        my_rom[2476] = 8'h8;
        my_rom[2477] = 8'h8;
        my_rom[2478] = 8'ha5;
        my_rom[2479] = 8'h5b;
        my_rom[2480] = 8'h53;
        my_rom[2481] = 8'h53;
        my_rom[2482] = 8'h53;
        my_rom[2483] = 8'h5b;
        my_rom[2484] = 8'h5b;
        my_rom[2485] = 8'h53;
        my_rom[2486] = 8'h53;
        my_rom[2487] = 8'h53;
        my_rom[2488] = 8'h53;
        my_rom[2489] = 8'h53;
        my_rom[2490] = 8'h53;
        my_rom[2491] = 8'h53;
        my_rom[2492] = 8'h53;
        my_rom[2493] = 8'h5b;
        my_rom[2494] = 8'h5b;
        my_rom[2495] = 8'h5b;
        my_rom[2496] = 8'h5b;
        my_rom[2497] = 8'h5b;
        my_rom[2498] = 8'h53;
        my_rom[2499] = 8'h53;
        my_rom[2500] = 8'h53;
        my_rom[2501] = 8'h53;
        my_rom[2502] = 8'h53;
        my_rom[2503] = 8'h53;
        my_rom[2504] = 8'h53;
        my_rom[2505] = 8'h4b;
        my_rom[2506] = 8'h49;
        my_rom[2507] = 8'h9;
        my_rom[2508] = 8'h9;
        my_rom[2509] = 8'h9;
        my_rom[2510] = 8'h9;
        my_rom[2511] = 8'h9;
        my_rom[2512] = 8'h9;
        my_rom[2513] = 8'h9;
        my_rom[2514] = 8'h9;
        my_rom[2515] = 8'h9;
        my_rom[2516] = 8'h9;
        my_rom[2517] = 8'hb;
        my_rom[2518] = 8'hb;
        my_rom[2519] = 8'h4b;
        my_rom[2520] = 8'h4b;
        my_rom[2521] = 8'h53;
        my_rom[2522] = 8'h53;
        my_rom[2523] = 8'h53;
        my_rom[2524] = 8'h8;
        my_rom[2525] = 8'h8;
        my_rom[2526] = 8'h8;
        my_rom[2527] = 8'h8;
        my_rom[2528] = 8'h8;
        my_rom[2529] = 8'h8;
        my_rom[2530] = 8'h8;
        my_rom[2531] = 8'ha;
        my_rom[2532] = 8'h8;
        my_rom[2533] = 8'h8;
        my_rom[2534] = 8'h8;
        my_rom[2535] = 8'h8;
        my_rom[2536] = 8'h8;
        my_rom[2537] = 8'hed;
        my_rom[2538] = 8'ha5;
        my_rom[2539] = 8'h9b;
        my_rom[2540] = 8'h9b;
        my_rom[2541] = 8'h9b;
        my_rom[2542] = 8'h9b;
        my_rom[2543] = 8'h5b;
        my_rom[2544] = 8'h9b;
        my_rom[2545] = 8'h9b;
        my_rom[2546] = 8'h9b;
        my_rom[2547] = 8'h9b;
        my_rom[2548] = 8'h9b;
        my_rom[2549] = 8'h9b;
        my_rom[2550] = 8'h9b;
        my_rom[2551] = 8'h9b;
        my_rom[2552] = 8'h9b;
        my_rom[2553] = 8'ha5;
        my_rom[2554] = 8'ha5;
        my_rom[2555] = 8'ha5;
        my_rom[2556] = 8'ha5;
        my_rom[2557] = 8'ha5;
        my_rom[2558] = 8'ha5;
        my_rom[2559] = 8'h9b;
        my_rom[2560] = 8'h9b;
        my_rom[2561] = 8'h5b;
        my_rom[2562] = 8'h5b;
        my_rom[2563] = 8'h53;
        my_rom[2564] = 8'h53;
        my_rom[2565] = 8'h53;
        my_rom[2566] = 8'h4b;
        my_rom[2567] = 8'h49;
        my_rom[2568] = 8'h49;
        my_rom[2569] = 8'h9;
        my_rom[2570] = 8'h9;
        my_rom[2571] = 8'h9;
        my_rom[2572] = 8'h9;
        my_rom[2573] = 8'h9;
        my_rom[2574] = 8'h9;
        my_rom[2575] = 8'h9;
        my_rom[2576] = 8'h9;
        my_rom[2577] = 8'h4b;
        my_rom[2578] = 8'h4b;
        my_rom[2579] = 8'h49;
        my_rom[2580] = 8'h49;
        my_rom[2581] = 8'h53;
        my_rom[2582] = 8'h53;
        my_rom[2583] = 8'h5b;
        my_rom[2584] = 8'h53;
        my_rom[2585] = 8'h8;
        my_rom[2586] = 8'h8;
        my_rom[2587] = 8'h8;
        my_rom[2588] = 8'h8;
        my_rom[2589] = 8'h8;
        my_rom[2590] = 8'h8;
        my_rom[2591] = 8'ha;
        my_rom[2592] = 8'h8;
        my_rom[2593] = 8'h8;
        my_rom[2594] = 8'h8;
        my_rom[2595] = 8'h8;
        my_rom[2596] = 8'hf7;
        my_rom[2597] = 8'had;
        my_rom[2598] = 8'h9b;
        my_rom[2599] = 8'h9b;
        my_rom[2600] = 8'h9b;
        my_rom[2601] = 8'h9b;
        my_rom[2602] = 8'h5b;
        my_rom[2603] = 8'h9b;
        my_rom[2604] = 8'h9b;
        my_rom[2605] = 8'h9b;
        my_rom[2606] = 8'h5b;
        my_rom[2607] = 8'h9b;
        my_rom[2608] = 8'ha3;
        my_rom[2609] = 8'ha5;
        my_rom[2610] = 8'ha5;
        my_rom[2611] = 8'had;
        my_rom[2612] = 8'hed;
        my_rom[2613] = 8'hed;
        my_rom[2614] = 8'hed;
        my_rom[2615] = 8'hed;
        my_rom[2616] = 8'hf7;
        my_rom[2617] = 8'hf7;
        my_rom[2618] = 8'hed;
        my_rom[2619] = 8'hed;
        my_rom[2620] = 8'had;
        my_rom[2621] = 8'ha5;
        my_rom[2622] = 8'ha3;
        my_rom[2623] = 8'h9b;
        my_rom[2624] = 8'h53;
        my_rom[2625] = 8'h51;
        my_rom[2626] = 8'h51;
        my_rom[2627] = 8'h4b;
        my_rom[2628] = 8'h49;
        my_rom[2629] = 8'h49;
        my_rom[2630] = 8'h49;
        my_rom[2631] = 8'h9;
        my_rom[2632] = 8'h9;
        my_rom[2633] = 8'h9;
        my_rom[2634] = 8'h9;
        my_rom[2635] = 8'h49;
        my_rom[2636] = 8'h49;
        my_rom[2637] = 8'h49;
        my_rom[2638] = 8'h49;
        my_rom[2639] = 8'h9;
        my_rom[2640] = 8'h9;
        my_rom[2641] = 8'h49;
        my_rom[2642] = 8'h49;
        my_rom[2643] = 8'h53;
        my_rom[2644] = 8'h5b;
        my_rom[2645] = 8'h8;
        my_rom[2646] = 8'h8;
        my_rom[2647] = 8'h8;
        my_rom[2648] = 8'h8;
        my_rom[2649] = 8'h8;
        my_rom[2650] = 8'h8;
        my_rom[2651] = 8'ha;
        my_rom[2652] = 8'h8;
        my_rom[2653] = 8'h8;
        my_rom[2654] = 8'h8;
        my_rom[2655] = 8'h8;
        my_rom[2656] = 8'hf7;
        my_rom[2657] = 8'ha5;
        my_rom[2658] = 8'h9b;
        my_rom[2659] = 8'h5b;
        my_rom[2660] = 8'h9b;
        my_rom[2661] = 8'h9b;
        my_rom[2662] = 8'h9b;
        my_rom[2663] = 8'h5b;
        my_rom[2664] = 8'h5b;
        my_rom[2665] = 8'h53;
        my_rom[2666] = 8'h5b;
        my_rom[2667] = 8'ha5;
        my_rom[2668] = 8'had;
        my_rom[2669] = 8'hed;
        my_rom[2670] = 8'hf7;
        my_rom[2671] = 8'hf7;
        my_rom[2672] = 8'hf7;
        my_rom[2673] = 8'hf7;
        my_rom[2674] = 8'hf7;
        my_rom[2675] = 8'hf7;
        my_rom[2676] = 8'hf7;
        my_rom[2677] = 8'hf7;
        my_rom[2678] = 8'hf7;
        my_rom[2679] = 8'hf7;
        my_rom[2680] = 8'hf7;
        my_rom[2681] = 8'hf7;
        my_rom[2682] = 8'hf7;
        my_rom[2683] = 8'hed;
        my_rom[2684] = 8'ha5;
        my_rom[2685] = 8'ha3;
        my_rom[2686] = 8'h5b;
        my_rom[2687] = 8'h53;
        my_rom[2688] = 8'h49;
        my_rom[2689] = 8'h49;
        my_rom[2690] = 8'h49;
        my_rom[2691] = 8'h49;
        my_rom[2692] = 8'h49;
        my_rom[2693] = 8'h49;
        my_rom[2694] = 8'h49;
        my_rom[2695] = 8'h49;
        my_rom[2696] = 8'h49;
        my_rom[2697] = 8'h49;
        my_rom[2698] = 8'h49;
        my_rom[2699] = 8'h49;
        my_rom[2700] = 8'h49;
        my_rom[2701] = 8'h49;
        my_rom[2702] = 8'h49;
        my_rom[2703] = 8'h53;
        my_rom[2704] = 8'h5b;
        my_rom[2705] = 8'h5b;
        my_rom[2706] = 8'h8;
        my_rom[2707] = 8'h8;
        my_rom[2708] = 8'h8;
        my_rom[2709] = 8'h8;
        my_rom[2710] = 8'h8;
        my_rom[2711] = 8'ha;
        my_rom[2712] = 8'h8;
        my_rom[2713] = 8'h8;
        my_rom[2714] = 8'h8;
        my_rom[2715] = 8'h8;
        my_rom[2716] = 8'ha5;
        my_rom[2717] = 8'h9b;
        my_rom[2718] = 8'h5b;
        my_rom[2719] = 8'h9b;
        my_rom[2720] = 8'h9b;
        my_rom[2721] = 8'h9b;
        my_rom[2722] = 8'h53;
        my_rom[2723] = 8'h5b;
        my_rom[2724] = 8'h9b;
        my_rom[2725] = 8'h53;
        my_rom[2726] = 8'ha3;
        my_rom[2727] = 8'hed;
        my_rom[2728] = 8'hf7;
        my_rom[2729] = 8'hf7;
        my_rom[2730] = 8'hf7;
        my_rom[2731] = 8'hf7;
        my_rom[2732] = 8'hf7;
        my_rom[2733] = 8'hf7;
        my_rom[2734] = 8'hf7;
        my_rom[2735] = 8'hf7;
        my_rom[2736] = 8'hf7;
        my_rom[2737] = 8'hf7;
        my_rom[2738] = 8'hf7;
        my_rom[2739] = 8'hf7;
        my_rom[2740] = 8'hf7;
        my_rom[2741] = 8'hf7;
        my_rom[2742] = 8'hf7;
        my_rom[2743] = 8'hf7;
        my_rom[2744] = 8'hf7;
        my_rom[2745] = 8'hed;
        my_rom[2746] = 8'hed;
        my_rom[2747] = 8'ha5;
        my_rom[2748] = 8'h9b;
        my_rom[2749] = 8'h9b;
        my_rom[2750] = 8'h53;
        my_rom[2751] = 8'h53;
        my_rom[2752] = 8'h53;
        my_rom[2753] = 8'h53;
        my_rom[2754] = 8'h53;
        my_rom[2755] = 8'h53;
        my_rom[2756] = 8'h51;
        my_rom[2757] = 8'h49;
        my_rom[2758] = 8'h49;
        my_rom[2759] = 8'h49;
        my_rom[2760] = 8'h49;
        my_rom[2761] = 8'h49;
        my_rom[2762] = 8'h51;
        my_rom[2763] = 8'h53;
        my_rom[2764] = 8'h5b;
        my_rom[2765] = 8'h5b;
        my_rom[2766] = 8'h8;
        my_rom[2767] = 8'h8;
        my_rom[2768] = 8'h8;
        my_rom[2769] = 8'h8;
        my_rom[2770] = 8'h8;
        my_rom[2771] = 8'ha;
        my_rom[2772] = 8'h8;
        my_rom[2773] = 8'h8;
        my_rom[2774] = 8'h8;
        my_rom[2775] = 8'h8;
        my_rom[2776] = 8'ha5;
        my_rom[2777] = 8'h5b;
        my_rom[2778] = 8'h9b;
        my_rom[2779] = 8'h9b;
        my_rom[2780] = 8'h5b;
        my_rom[2781] = 8'h53;
        my_rom[2782] = 8'h53;
        my_rom[2783] = 8'h9b;
        my_rom[2784] = 8'h53;
        my_rom[2785] = 8'h5b;
        my_rom[2786] = 8'had;
        my_rom[2787] = 8'hf7;
        my_rom[2788] = 8'hf7;
        my_rom[2789] = 8'hf7;
        my_rom[2790] = 8'hf7;
        my_rom[2791] = 8'hf7;
        my_rom[2792] = 8'hf7;
        my_rom[2793] = 8'hf7;
        my_rom[2794] = 8'hf7;
        my_rom[2795] = 8'hf7;
        my_rom[2796] = 8'hf7;
        my_rom[2797] = 8'hf7;
        my_rom[2798] = 8'hf7;
        my_rom[2799] = 8'hf7;
        my_rom[2800] = 8'hf7;
        my_rom[2801] = 8'hf7;
        my_rom[2802] = 8'hf7;
        my_rom[2803] = 8'hf7;
        my_rom[2804] = 8'hf7;
        my_rom[2805] = 8'hf7;
        my_rom[2806] = 8'hf7;
        my_rom[2807] = 8'hef;
        my_rom[2808] = 8'hed;
        my_rom[2809] = 8'had;
        my_rom[2810] = 8'ha5;
        my_rom[2811] = 8'ha5;
        my_rom[2812] = 8'ha5;
        my_rom[2813] = 8'ha5;
        my_rom[2814] = 8'h9d;
        my_rom[2815] = 8'h9b;
        my_rom[2816] = 8'h9b;
        my_rom[2817] = 8'h53;
        my_rom[2818] = 8'h49;
        my_rom[2819] = 8'h49;
        my_rom[2820] = 8'h49;
        my_rom[2821] = 8'h9;
        my_rom[2822] = 8'h53;
        my_rom[2823] = 8'h53;
        my_rom[2824] = 8'h53;
        my_rom[2825] = 8'ha3;
        my_rom[2826] = 8'ha3;
        my_rom[2827] = 8'h8;
        my_rom[2828] = 8'h8;
        my_rom[2829] = 8'h8;
        my_rom[2830] = 8'h8;
        my_rom[2831] = 8'ha;
        my_rom[2832] = 8'h8;
        my_rom[2833] = 8'h8;
        my_rom[2834] = 8'h8;
        my_rom[2835] = 8'hf7;
        my_rom[2836] = 8'ha5;
        my_rom[2837] = 8'h53;
        my_rom[2838] = 8'h9b;
        my_rom[2839] = 8'h9b;
        my_rom[2840] = 8'h53;
        my_rom[2841] = 8'h53;
        my_rom[2842] = 8'h53;
        my_rom[2843] = 8'h9b;
        my_rom[2844] = 8'h53;
        my_rom[2845] = 8'h9b;
        my_rom[2846] = 8'hed;
        my_rom[2847] = 8'hf7;
        my_rom[2848] = 8'hf7;
        my_rom[2849] = 8'hf7;
        my_rom[2850] = 8'hf7;
        my_rom[2851] = 8'hf7;
        my_rom[2852] = 8'hf7;
        my_rom[2853] = 8'hf7;
        my_rom[2854] = 8'hf7;
        my_rom[2855] = 8'hf7;
        my_rom[2856] = 8'hf7;
        my_rom[2857] = 8'hf7;
        my_rom[2858] = 8'hf7;
        my_rom[2859] = 8'hf7;
        my_rom[2860] = 8'hf7;
        my_rom[2861] = 8'hf7;
        my_rom[2862] = 8'hf7;
        my_rom[2863] = 8'hf7;
        my_rom[2864] = 8'hf7;
        my_rom[2865] = 8'hf7;
        my_rom[2866] = 8'hf7;
        my_rom[2867] = 8'hf7;
        my_rom[2868] = 8'hf7;
        my_rom[2869] = 8'hef;
        my_rom[2870] = 8'hef;
        my_rom[2871] = 8'haf;
        my_rom[2872] = 8'had;
        my_rom[2873] = 8'had;
        my_rom[2874] = 8'had;
        my_rom[2875] = 8'had;
        my_rom[2876] = 8'had;
        my_rom[2877] = 8'ha5;
        my_rom[2878] = 8'h9b;
        my_rom[2879] = 8'h49;
        my_rom[2880] = 8'h9;
        my_rom[2881] = 8'h9;
        my_rom[2882] = 8'h9;
        my_rom[2883] = 8'h53;
        my_rom[2884] = 8'h53;
        my_rom[2885] = 8'h9b;
        my_rom[2886] = 8'ha3;
        my_rom[2887] = 8'h8;
        my_rom[2888] = 8'h8;
        my_rom[2889] = 8'h8;
        my_rom[2890] = 8'h8;
        my_rom[2891] = 8'ha;
        my_rom[2892] = 8'h8;
        my_rom[2893] = 8'h8;
        my_rom[2894] = 8'h8;
        my_rom[2895] = 8'hf7;
        my_rom[2896] = 8'h9b;
        my_rom[2897] = 8'h53;
        my_rom[2898] = 8'h9b;
        my_rom[2899] = 8'h9b;
        my_rom[2900] = 8'h53;
        my_rom[2901] = 8'h53;
        my_rom[2902] = 8'h5b;
        my_rom[2903] = 8'h5b;
        my_rom[2904] = 8'h5b;
        my_rom[2905] = 8'had;
        my_rom[2906] = 8'hf7;
        my_rom[2907] = 8'hf7;
        my_rom[2908] = 8'hf7;
        my_rom[2909] = 8'hf7;
        my_rom[2910] = 8'hf7;
        my_rom[2911] = 8'hf7;
        my_rom[2912] = 8'hff;
        my_rom[2913] = 8'hff;
        my_rom[2914] = 8'hff;
        my_rom[2915] = 8'hf7;
        my_rom[2916] = 8'hf7;
        my_rom[2917] = 8'hf7;
        my_rom[2918] = 8'hf7;
        my_rom[2919] = 8'hf7;
        my_rom[2920] = 8'hf7;
        my_rom[2921] = 8'hf7;
        my_rom[2922] = 8'hf7;
        my_rom[2923] = 8'hf7;
        my_rom[2924] = 8'hf7;
        my_rom[2925] = 8'hf7;
        my_rom[2926] = 8'hf7;
        my_rom[2927] = 8'hf7;
        my_rom[2928] = 8'hf7;
        my_rom[2929] = 8'hf7;
        my_rom[2930] = 8'hf7;
        my_rom[2931] = 8'hf7;
        my_rom[2932] = 8'hf7;
        my_rom[2933] = 8'haf;
        my_rom[2934] = 8'haf;
        my_rom[2935] = 8'haf;
        my_rom[2936] = 8'haf;
        my_rom[2937] = 8'haf;
        my_rom[2938] = 8'had;
        my_rom[2939] = 8'ha5;
        my_rom[2940] = 8'h49;
        my_rom[2941] = 8'h49;
        my_rom[2942] = 8'h49;
        my_rom[2943] = 8'h4b;
        my_rom[2944] = 8'h53;
        my_rom[2945] = 8'h5b;
        my_rom[2946] = 8'ha3;
        my_rom[2947] = 8'h8;
        my_rom[2948] = 8'h8;
        my_rom[2949] = 8'h8;
        my_rom[2950] = 8'h8;
        my_rom[2951] = 8'ha;
        my_rom[2952] = 8'h8;
        my_rom[2953] = 8'h8;
        my_rom[2954] = 8'h8;
        my_rom[2955] = 8'had;
        my_rom[2956] = 8'h5b;
        my_rom[2957] = 8'h5b;
        my_rom[2958] = 8'ha3;
        my_rom[2959] = 8'h9b;
        my_rom[2960] = 8'h53;
        my_rom[2961] = 8'h9b;
        my_rom[2962] = 8'h9b;
        my_rom[2963] = 8'h5b;
        my_rom[2964] = 8'ha5;
        my_rom[2965] = 8'hed;
        my_rom[2966] = 8'hf7;
        my_rom[2967] = 8'hf7;
        my_rom[2968] = 8'hf7;
        my_rom[2969] = 8'hf7;
        my_rom[2970] = 8'hf7;
        my_rom[2971] = 8'hff;
        my_rom[2972] = 8'hff;
        my_rom[2973] = 8'hff;
        my_rom[2974] = 8'hff;
        my_rom[2975] = 8'hff;
        my_rom[2976] = 8'hf7;
        my_rom[2977] = 8'hf7;
        my_rom[2978] = 8'hf7;
        my_rom[2979] = 8'hf7;
        my_rom[2980] = 8'hf7;
        my_rom[2981] = 8'hf7;
        my_rom[2982] = 8'hf7;
        my_rom[2983] = 8'hf7;
        my_rom[2984] = 8'hf7;
        my_rom[2985] = 8'hf7;
        my_rom[2986] = 8'hf7;
        my_rom[2987] = 8'hf7;
        my_rom[2988] = 8'hf7;
        my_rom[2989] = 8'hf7;
        my_rom[2990] = 8'hf7;
        my_rom[2991] = 8'hf7;
        my_rom[2992] = 8'hf7;
        my_rom[2993] = 8'hef;
        my_rom[2994] = 8'hef;
        my_rom[2995] = 8'haf;
        my_rom[2996] = 8'haf;
        my_rom[2997] = 8'haf;
        my_rom[2998] = 8'haf;
        my_rom[2999] = 8'haf;
        my_rom[3000] = 8'h9d;
        my_rom[3001] = 8'h53;
        my_rom[3002] = 8'h49;
        my_rom[3003] = 8'h4b;
        my_rom[3004] = 8'h53;
        my_rom[3005] = 8'h53;
        my_rom[3006] = 8'ha3;
        my_rom[3007] = 8'ha3;
        my_rom[3008] = 8'h8;
        my_rom[3009] = 8'h8;
        my_rom[3010] = 8'h8;
        my_rom[3011] = 8'ha;
        my_rom[3012] = 8'h8;
        my_rom[3013] = 8'h8;
        my_rom[3014] = 8'h8;
        my_rom[3015] = 8'ha5;
        my_rom[3016] = 8'h53;
        my_rom[3017] = 8'h5b;
        my_rom[3018] = 8'h9b;
        my_rom[3019] = 8'h9b;
        my_rom[3020] = 8'h5b;
        my_rom[3021] = 8'h9b;
        my_rom[3022] = 8'h5b;
        my_rom[3023] = 8'h5b;
        my_rom[3024] = 8'ha5;
        my_rom[3025] = 8'hed;
        my_rom[3026] = 8'hf7;
        my_rom[3027] = 8'hf7;
        my_rom[3028] = 8'hf7;
        my_rom[3029] = 8'hf7;
        my_rom[3030] = 8'hff;
        my_rom[3031] = 8'hff;
        my_rom[3032] = 8'hff;
        my_rom[3033] = 8'hff;
        my_rom[3034] = 8'hff;
        my_rom[3035] = 8'hf7;
        my_rom[3036] = 8'hf7;
        my_rom[3037] = 8'hf7;
        my_rom[3038] = 8'hf7;
        my_rom[3039] = 8'hf7;
        my_rom[3040] = 8'hf7;
        my_rom[3041] = 8'hf7;
        my_rom[3042] = 8'hf7;
        my_rom[3043] = 8'hf7;
        my_rom[3044] = 8'hf7;
        my_rom[3045] = 8'hf7;
        my_rom[3046] = 8'hf7;
        my_rom[3047] = 8'hf7;
        my_rom[3048] = 8'hf7;
        my_rom[3049] = 8'hf7;
        my_rom[3050] = 8'hf7;
        my_rom[3051] = 8'hf7;
        my_rom[3052] = 8'hef;
        my_rom[3053] = 8'hef;
        my_rom[3054] = 8'hef;
        my_rom[3055] = 8'hef;
        my_rom[3056] = 8'haf;
        my_rom[3057] = 8'hef;
        my_rom[3058] = 8'haf;
        my_rom[3059] = 8'haf;
        my_rom[3060] = 8'ha5;
        my_rom[3061] = 8'h5b;
        my_rom[3062] = 8'h53;
        my_rom[3063] = 8'h53;
        my_rom[3064] = 8'h53;
        my_rom[3065] = 8'h53;
        my_rom[3066] = 8'ha3;
        my_rom[3067] = 8'ha3;
        my_rom[3068] = 8'h8;
        my_rom[3069] = 8'h8;
        my_rom[3070] = 8'h8;
        my_rom[3071] = 8'ha;
        my_rom[3072] = 8'h8;
        my_rom[3073] = 8'h8;
        my_rom[3074] = 8'hf7;
        my_rom[3075] = 8'h9b;
        my_rom[3076] = 8'h53;
        my_rom[3077] = 8'h5b;
        my_rom[3078] = 8'h9b;
        my_rom[3079] = 8'h5b;
        my_rom[3080] = 8'h9b;
        my_rom[3081] = 8'ha3;
        my_rom[3082] = 8'h53;
        my_rom[3083] = 8'h5b;
        my_rom[3084] = 8'ha5;
        my_rom[3085] = 8'hed;
        my_rom[3086] = 8'hf7;
        my_rom[3087] = 8'hf7;
        my_rom[3088] = 8'hf7;
        my_rom[3089] = 8'hff;
        my_rom[3090] = 8'hff;
        my_rom[3091] = 8'hf7;
        my_rom[3092] = 8'hff;
        my_rom[3093] = 8'hff;
        my_rom[3094] = 8'hf7;
        my_rom[3095] = 8'hf7;
        my_rom[3096] = 8'hf7;
        my_rom[3097] = 8'hf7;
        my_rom[3098] = 8'hf7;
        my_rom[3099] = 8'hf7;
        my_rom[3100] = 8'hf7;
        my_rom[3101] = 8'hf7;
        my_rom[3102] = 8'hf7;
        my_rom[3103] = 8'hf7;
        my_rom[3104] = 8'hf7;
        my_rom[3105] = 8'hf7;
        my_rom[3106] = 8'hf7;
        my_rom[3107] = 8'hf7;
        my_rom[3108] = 8'hf7;
        my_rom[3109] = 8'hf7;
        my_rom[3110] = 8'hf7;
        my_rom[3111] = 8'hef;
        my_rom[3112] = 8'hef;
        my_rom[3113] = 8'hef;
        my_rom[3114] = 8'hef;
        my_rom[3115] = 8'hef;
        my_rom[3116] = 8'hef;
        my_rom[3117] = 8'haf;
        my_rom[3118] = 8'haf;
        my_rom[3119] = 8'haf;
        my_rom[3120] = 8'had;
        my_rom[3121] = 8'h5d;
        my_rom[3122] = 8'h53;
        my_rom[3123] = 8'h53;
        my_rom[3124] = 8'h53;
        my_rom[3125] = 8'h53;
        my_rom[3126] = 8'h5b;
        my_rom[3127] = 8'had;
        my_rom[3128] = 8'h8;
        my_rom[3129] = 8'h8;
        my_rom[3130] = 8'h8;
        my_rom[3131] = 8'ha;
        my_rom[3132] = 8'h8;
        my_rom[3133] = 8'h8;
        my_rom[3134] = 8'hf7;
        my_rom[3135] = 8'h5b;
        my_rom[3136] = 8'h53;
        my_rom[3137] = 8'h9b;
        my_rom[3138] = 8'h9b;
        my_rom[3139] = 8'h5b;
        my_rom[3140] = 8'h9b;
        my_rom[3141] = 8'h5b;
        my_rom[3142] = 8'h53;
        my_rom[3143] = 8'h5b;
        my_rom[3144] = 8'had;
        my_rom[3145] = 8'hed;
        my_rom[3146] = 8'hf7;
        my_rom[3147] = 8'hf7;
        my_rom[3148] = 8'hf7;
        my_rom[3149] = 8'hf7;
        my_rom[3150] = 8'hf7;
        my_rom[3151] = 8'hf7;
        my_rom[3152] = 8'hf7;
        my_rom[3153] = 8'hf7;
        my_rom[3154] = 8'hf7;
        my_rom[3155] = 8'hf7;
        my_rom[3156] = 8'hf7;
        my_rom[3157] = 8'hf7;
        my_rom[3158] = 8'hf7;
        my_rom[3159] = 8'hf7;
        my_rom[3160] = 8'hf7;
        my_rom[3161] = 8'hf7;
        my_rom[3162] = 8'hf7;
        my_rom[3163] = 8'hf7;
        my_rom[3164] = 8'hf7;
        my_rom[3165] = 8'hf7;
        my_rom[3166] = 8'hf7;
        my_rom[3167] = 8'hf7;
        my_rom[3168] = 8'hf7;
        my_rom[3169] = 8'hef;
        my_rom[3170] = 8'hef;
        my_rom[3171] = 8'hef;
        my_rom[3172] = 8'hef;
        my_rom[3173] = 8'hef;
        my_rom[3174] = 8'hef;
        my_rom[3175] = 8'haf;
        my_rom[3176] = 8'haf;
        my_rom[3177] = 8'haf;
        my_rom[3178] = 8'hef;
        my_rom[3179] = 8'hef;
        my_rom[3180] = 8'had;
        my_rom[3181] = 8'ha5;
        my_rom[3182] = 8'h53;
        my_rom[3183] = 8'h4b;
        my_rom[3184] = 8'h53;
        my_rom[3185] = 8'h53;
        my_rom[3186] = 8'h53;
        my_rom[3187] = 8'had;
        my_rom[3188] = 8'h8;
        my_rom[3189] = 8'h8;
        my_rom[3190] = 8'h8;
        my_rom[3191] = 8'ha;
        my_rom[3192] = 8'h8;
        my_rom[3193] = 8'h8;
        my_rom[3194] = 8'hed;
        my_rom[3195] = 8'h5b;
        my_rom[3196] = 8'h5b;
        my_rom[3197] = 8'h9b;
        my_rom[3198] = 8'h9b;
        my_rom[3199] = 8'h53;
        my_rom[3200] = 8'h53;
        my_rom[3201] = 8'h53;
        my_rom[3202] = 8'h53;
        my_rom[3203] = 8'h9b;
        my_rom[3204] = 8'had;
        my_rom[3205] = 8'hed;
        my_rom[3206] = 8'hf7;
        my_rom[3207] = 8'hf7;
        my_rom[3208] = 8'hf7;
        my_rom[3209] = 8'hf7;
        my_rom[3210] = 8'hf7;
        my_rom[3211] = 8'hf7;
        my_rom[3212] = 8'hf7;
        my_rom[3213] = 8'hf7;
        my_rom[3214] = 8'hf7;
        my_rom[3215] = 8'hf7;
        my_rom[3216] = 8'hf7;
        my_rom[3217] = 8'hf7;
        my_rom[3218] = 8'hf7;
        my_rom[3219] = 8'hf7;
        my_rom[3220] = 8'hf7;
        my_rom[3221] = 8'hf7;
        my_rom[3222] = 8'hf7;
        my_rom[3223] = 8'hf7;
        my_rom[3224] = 8'hf7;
        my_rom[3225] = 8'hf7;
        my_rom[3226] = 8'hf7;
        my_rom[3227] = 8'hf7;
        my_rom[3228] = 8'hef;
        my_rom[3229] = 8'hef;
        my_rom[3230] = 8'hef;
        my_rom[3231] = 8'hef;
        my_rom[3232] = 8'hef;
        my_rom[3233] = 8'hef;
        my_rom[3234] = 8'haf;
        my_rom[3235] = 8'haf;
        my_rom[3236] = 8'haf;
        my_rom[3237] = 8'haf;
        my_rom[3238] = 8'haf;
        my_rom[3239] = 8'hef;
        my_rom[3240] = 8'had;
        my_rom[3241] = 8'ha5;
        my_rom[3242] = 8'h53;
        my_rom[3243] = 8'h4b;
        my_rom[3244] = 8'h53;
        my_rom[3245] = 8'h53;
        my_rom[3246] = 8'h53;
        my_rom[3247] = 8'had;
        my_rom[3248] = 8'h8;
        my_rom[3249] = 8'h8;
        my_rom[3250] = 8'h8;
        my_rom[3251] = 8'ha;
        my_rom[3252] = 8'h8;
        my_rom[3253] = 8'h8;
        my_rom[3254] = 8'had;
        my_rom[3255] = 8'h5b;
        my_rom[3256] = 8'h5b;
        my_rom[3257] = 8'h9b;
        my_rom[3258] = 8'h53;
        my_rom[3259] = 8'h53;
        my_rom[3260] = 8'h53;
        my_rom[3261] = 8'h53;
        my_rom[3262] = 8'h53;
        my_rom[3263] = 8'ha5;
        my_rom[3264] = 8'had;
        my_rom[3265] = 8'hed;
        my_rom[3266] = 8'hf7;
        my_rom[3267] = 8'hf7;
        my_rom[3268] = 8'hf7;
        my_rom[3269] = 8'hf7;
        my_rom[3270] = 8'hf7;
        my_rom[3271] = 8'hf7;
        my_rom[3272] = 8'hf7;
        my_rom[3273] = 8'hf7;
        my_rom[3274] = 8'hf7;
        my_rom[3275] = 8'hf7;
        my_rom[3276] = 8'hf7;
        my_rom[3277] = 8'hf7;
        my_rom[3278] = 8'hf7;
        my_rom[3279] = 8'hf7;
        my_rom[3280] = 8'hf7;
        my_rom[3281] = 8'hf7;
        my_rom[3282] = 8'hf7;
        my_rom[3283] = 8'hf7;
        my_rom[3284] = 8'hf7;
        my_rom[3285] = 8'hf7;
        my_rom[3286] = 8'hf7;
        my_rom[3287] = 8'hf7;
        my_rom[3288] = 8'hef;
        my_rom[3289] = 8'hef;
        my_rom[3290] = 8'hef;
        my_rom[3291] = 8'hef;
        my_rom[3292] = 8'hef;
        my_rom[3293] = 8'hef;
        my_rom[3294] = 8'haf;
        my_rom[3295] = 8'haf;
        my_rom[3296] = 8'haf;
        my_rom[3297] = 8'haf;
        my_rom[3298] = 8'haf;
        my_rom[3299] = 8'hef;
        my_rom[3300] = 8'had;
        my_rom[3301] = 8'ha5;
        my_rom[3302] = 8'h5b;
        my_rom[3303] = 8'h53;
        my_rom[3304] = 8'h49;
        my_rom[3305] = 8'h51;
        my_rom[3306] = 8'h53;
        my_rom[3307] = 8'had;
        my_rom[3308] = 8'hed;
        my_rom[3309] = 8'h8;
        my_rom[3310] = 8'h8;
        my_rom[3311] = 8'ha;
        my_rom[3312] = 8'h8;
        my_rom[3313] = 8'h8;
        my_rom[3314] = 8'ha5;
        my_rom[3315] = 8'h53;
        my_rom[3316] = 8'h53;
        my_rom[3317] = 8'h5b;
        my_rom[3318] = 8'h53;
        my_rom[3319] = 8'h53;
        my_rom[3320] = 8'h53;
        my_rom[3321] = 8'h4b;
        my_rom[3322] = 8'h5b;
        my_rom[3323] = 8'ha5;
        my_rom[3324] = 8'had;
        my_rom[3325] = 8'hed;
        my_rom[3326] = 8'hf7;
        my_rom[3327] = 8'hf7;
        my_rom[3328] = 8'hf7;
        my_rom[3329] = 8'hf7;
        my_rom[3330] = 8'hf7;
        my_rom[3331] = 8'hf7;
        my_rom[3332] = 8'hf7;
        my_rom[3333] = 8'hf7;
        my_rom[3334] = 8'hf7;
        my_rom[3335] = 8'hf7;
        my_rom[3336] = 8'hf7;
        my_rom[3337] = 8'hf7;
        my_rom[3338] = 8'hf7;
        my_rom[3339] = 8'hf7;
        my_rom[3340] = 8'hf7;
        my_rom[3341] = 8'hf7;
        my_rom[3342] = 8'hf7;
        my_rom[3343] = 8'hf7;
        my_rom[3344] = 8'hf7;
        my_rom[3345] = 8'hf7;
        my_rom[3346] = 8'hf7;
        my_rom[3347] = 8'hf7;
        my_rom[3348] = 8'hf7;
        my_rom[3349] = 8'hf7;
        my_rom[3350] = 8'hf7;
        my_rom[3351] = 8'hf7;
        my_rom[3352] = 8'hef;
        my_rom[3353] = 8'hef;
        my_rom[3354] = 8'haf;
        my_rom[3355] = 8'had;
        my_rom[3356] = 8'had;
        my_rom[3357] = 8'had;
        my_rom[3358] = 8'haf;
        my_rom[3359] = 8'hef;
        my_rom[3360] = 8'hed;
        my_rom[3361] = 8'ha5;
        my_rom[3362] = 8'h5b;
        my_rom[3363] = 8'h53;
        my_rom[3364] = 8'h49;
        my_rom[3365] = 8'h49;
        my_rom[3366] = 8'h53;
        my_rom[3367] = 8'had;
        my_rom[3368] = 8'hed;
        my_rom[3369] = 8'h8;
        my_rom[3370] = 8'h8;
        my_rom[3371] = 8'ha;
        my_rom[3372] = 8'h8;
        my_rom[3373] = 8'h8;
        my_rom[3374] = 8'ha5;
        my_rom[3375] = 8'h53;
        my_rom[3376] = 8'h53;
        my_rom[3377] = 8'h5b;
        my_rom[3378] = 8'h53;
        my_rom[3379] = 8'h53;
        my_rom[3380] = 8'h49;
        my_rom[3381] = 8'h53;
        my_rom[3382] = 8'h9b;
        my_rom[3383] = 8'ha5;
        my_rom[3384] = 8'ha5;
        my_rom[3385] = 8'hed;
        my_rom[3386] = 8'hf7;
        my_rom[3387] = 8'hf7;
        my_rom[3388] = 8'hf7;
        my_rom[3389] = 8'hf7;
        my_rom[3390] = 8'hf7;
        my_rom[3391] = 8'hf7;
        my_rom[3392] = 8'hf7;
        my_rom[3393] = 8'hf7;
        my_rom[3394] = 8'hf7;
        my_rom[3395] = 8'hf7;
        my_rom[3396] = 8'hf7;
        my_rom[3397] = 8'hf7;
        my_rom[3398] = 8'hf7;
        my_rom[3399] = 8'hf7;
        my_rom[3400] = 8'hf7;
        my_rom[3401] = 8'hf7;
        my_rom[3402] = 8'hf7;
        my_rom[3403] = 8'hf7;
        my_rom[3404] = 8'hf7;
        my_rom[3405] = 8'hf7;
        my_rom[3406] = 8'hf7;
        my_rom[3407] = 8'hf7;
        my_rom[3408] = 8'hf7;
        my_rom[3409] = 8'hf7;
        my_rom[3410] = 8'hf7;
        my_rom[3411] = 8'hf7;
        my_rom[3412] = 8'hf7;
        my_rom[3413] = 8'hef;
        my_rom[3414] = 8'hef;
        my_rom[3415] = 8'haf;
        my_rom[3416] = 8'haf;
        my_rom[3417] = 8'haf;
        my_rom[3418] = 8'haf;
        my_rom[3419] = 8'hef;
        my_rom[3420] = 8'had;
        my_rom[3421] = 8'had;
        my_rom[3422] = 8'h9b;
        my_rom[3423] = 8'h53;
        my_rom[3424] = 8'h49;
        my_rom[3425] = 8'h49;
        my_rom[3426] = 8'h49;
        my_rom[3427] = 8'ha3;
        my_rom[3428] = 8'hed;
        my_rom[3429] = 8'h8;
        my_rom[3430] = 8'h8;
        my_rom[3431] = 8'ha;
        my_rom[3432] = 8'h8;
        my_rom[3433] = 8'h8;
        my_rom[3434] = 8'ha5;
        my_rom[3435] = 8'h53;
        my_rom[3436] = 8'h53;
        my_rom[3437] = 8'h53;
        my_rom[3438] = 8'h53;
        my_rom[3439] = 8'h53;
        my_rom[3440] = 8'h53;
        my_rom[3441] = 8'h53;
        my_rom[3442] = 8'h5b;
        my_rom[3443] = 8'ha5;
        my_rom[3444] = 8'ha5;
        my_rom[3445] = 8'had;
        my_rom[3446] = 8'hf7;
        my_rom[3447] = 8'hf7;
        my_rom[3448] = 8'hf7;
        my_rom[3449] = 8'hf7;
        my_rom[3450] = 8'hf7;
        my_rom[3451] = 8'hf7;
        my_rom[3452] = 8'hf7;
        my_rom[3453] = 8'hf7;
        my_rom[3454] = 8'hf7;
        my_rom[3455] = 8'hf7;
        my_rom[3456] = 8'hf7;
        my_rom[3457] = 8'hf7;
        my_rom[3458] = 8'hf7;
        my_rom[3459] = 8'hf7;
        my_rom[3460] = 8'hf7;
        my_rom[3461] = 8'hf7;
        my_rom[3462] = 8'hf7;
        my_rom[3463] = 8'hf7;
        my_rom[3464] = 8'hf7;
        my_rom[3465] = 8'hf7;
        my_rom[3466] = 8'hf7;
        my_rom[3467] = 8'hf7;
        my_rom[3468] = 8'hf7;
        my_rom[3469] = 8'hf7;
        my_rom[3470] = 8'hf7;
        my_rom[3471] = 8'hf7;
        my_rom[3472] = 8'hf7;
        my_rom[3473] = 8'hf7;
        my_rom[3474] = 8'hef;
        my_rom[3475] = 8'haf;
        my_rom[3476] = 8'haf;
        my_rom[3477] = 8'haf;
        my_rom[3478] = 8'haf;
        my_rom[3479] = 8'hef;
        my_rom[3480] = 8'had;
        my_rom[3481] = 8'had;
        my_rom[3482] = 8'h9d;
        my_rom[3483] = 8'h53;
        my_rom[3484] = 8'h49;
        my_rom[3485] = 8'h49;
        my_rom[3486] = 8'h49;
        my_rom[3487] = 8'ha3;
        my_rom[3488] = 8'hed;
        my_rom[3489] = 8'h8;
        my_rom[3490] = 8'h8;
        my_rom[3491] = 8'ha;
        my_rom[3492] = 8'h8;
        my_rom[3493] = 8'h8;
        my_rom[3494] = 8'ha5;
        my_rom[3495] = 8'h53;
        my_rom[3496] = 8'h53;
        my_rom[3497] = 8'h5b;
        my_rom[3498] = 8'h53;
        my_rom[3499] = 8'h53;
        my_rom[3500] = 8'h53;
        my_rom[3501] = 8'h53;
        my_rom[3502] = 8'h5b;
        my_rom[3503] = 8'h9b;
        my_rom[3504] = 8'ha5;
        my_rom[3505] = 8'hed;
        my_rom[3506] = 8'hf7;
        my_rom[3507] = 8'hf7;
        my_rom[3508] = 8'hf7;
        my_rom[3509] = 8'hf7;
        my_rom[3510] = 8'hf7;
        my_rom[3511] = 8'hf7;
        my_rom[3512] = 8'hf7;
        my_rom[3513] = 8'hf7;
        my_rom[3514] = 8'hf7;
        my_rom[3515] = 8'hf7;
        my_rom[3516] = 8'hf7;
        my_rom[3517] = 8'hf7;
        my_rom[3518] = 8'hf7;
        my_rom[3519] = 8'hf7;
        my_rom[3520] = 8'hf7;
        my_rom[3521] = 8'hf7;
        my_rom[3522] = 8'hf7;
        my_rom[3523] = 8'hf7;
        my_rom[3524] = 8'hf7;
        my_rom[3525] = 8'hf7;
        my_rom[3526] = 8'hf7;
        my_rom[3527] = 8'hf7;
        my_rom[3528] = 8'hf7;
        my_rom[3529] = 8'hf7;
        my_rom[3530] = 8'hf7;
        my_rom[3531] = 8'hf7;
        my_rom[3532] = 8'hf7;
        my_rom[3533] = 8'hf7;
        my_rom[3534] = 8'hf7;
        my_rom[3535] = 8'hef;
        my_rom[3536] = 8'hef;
        my_rom[3537] = 8'haf;
        my_rom[3538] = 8'haf;
        my_rom[3539] = 8'haf;
        my_rom[3540] = 8'had;
        my_rom[3541] = 8'had;
        my_rom[3542] = 8'ha5;
        my_rom[3543] = 8'h53;
        my_rom[3544] = 8'h49;
        my_rom[3545] = 8'h49;
        my_rom[3546] = 8'h49;
        my_rom[3547] = 8'h9b;
        my_rom[3548] = 8'had;
        my_rom[3549] = 8'h8;
        my_rom[3550] = 8'h8;
        my_rom[3551] = 8'ha;
        my_rom[3552] = 8'h8;
        my_rom[3553] = 8'h8;
        my_rom[3554] = 8'ha5;
        my_rom[3555] = 8'h53;
        my_rom[3556] = 8'h53;
        my_rom[3557] = 8'h53;
        my_rom[3558] = 8'h53;
        my_rom[3559] = 8'h53;
        my_rom[3560] = 8'h53;
        my_rom[3561] = 8'h53;
        my_rom[3562] = 8'h53;
        my_rom[3563] = 8'h5b;
        my_rom[3564] = 8'ha5;
        my_rom[3565] = 8'hed;
        my_rom[3566] = 8'hf7;
        my_rom[3567] = 8'hf7;
        my_rom[3568] = 8'hf7;
        my_rom[3569] = 8'hf7;
        my_rom[3570] = 8'hf7;
        my_rom[3571] = 8'hf7;
        my_rom[3572] = 8'hf7;
        my_rom[3573] = 8'hf7;
        my_rom[3574] = 8'hf7;
        my_rom[3575] = 8'hf7;
        my_rom[3576] = 8'hf7;
        my_rom[3577] = 8'hf7;
        my_rom[3578] = 8'hf7;
        my_rom[3579] = 8'hf7;
        my_rom[3580] = 8'hf7;
        my_rom[3581] = 8'hf7;
        my_rom[3582] = 8'hf7;
        my_rom[3583] = 8'hf7;
        my_rom[3584] = 8'hf7;
        my_rom[3585] = 8'hf7;
        my_rom[3586] = 8'hf7;
        my_rom[3587] = 8'hf7;
        my_rom[3588] = 8'hf7;
        my_rom[3589] = 8'hf7;
        my_rom[3590] = 8'hf7;
        my_rom[3591] = 8'hf7;
        my_rom[3592] = 8'hef;
        my_rom[3593] = 8'hef;
        my_rom[3594] = 8'haf;
        my_rom[3595] = 8'haf;
        my_rom[3596] = 8'haf;
        my_rom[3597] = 8'haf;
        my_rom[3598] = 8'haf;
        my_rom[3599] = 8'haf;
        my_rom[3600] = 8'haf;
        my_rom[3601] = 8'had;
        my_rom[3602] = 8'ha5;
        my_rom[3603] = 8'h53;
        my_rom[3604] = 8'h49;
        my_rom[3605] = 8'h49;
        my_rom[3606] = 8'h49;
        my_rom[3607] = 8'h5b;
        my_rom[3608] = 8'had;
        my_rom[3609] = 8'h8;
        my_rom[3610] = 8'h8;
        my_rom[3611] = 8'ha;
        my_rom[3612] = 8'h8;
        my_rom[3613] = 8'h8;
        my_rom[3614] = 8'ha5;
        my_rom[3615] = 8'h53;
        my_rom[3616] = 8'h53;
        my_rom[3617] = 8'h53;
        my_rom[3618] = 8'h53;
        my_rom[3619] = 8'h53;
        my_rom[3620] = 8'h53;
        my_rom[3621] = 8'h53;
        my_rom[3622] = 8'h53;
        my_rom[3623] = 8'h53;
        my_rom[3624] = 8'ha5;
        my_rom[3625] = 8'hed;
        my_rom[3626] = 8'hf7;
        my_rom[3627] = 8'hf7;
        my_rom[3628] = 8'hf7;
        my_rom[3629] = 8'hf7;
        my_rom[3630] = 8'hf7;
        my_rom[3631] = 8'hf7;
        my_rom[3632] = 8'had;
        my_rom[3633] = 8'ha5;
        my_rom[3634] = 8'ha5;
        my_rom[3635] = 8'ha5;
        my_rom[3636] = 8'ha5;
        my_rom[3637] = 8'ha5;
        my_rom[3638] = 8'ha5;
        my_rom[3639] = 8'ha5;
        my_rom[3640] = 8'had;
        my_rom[3641] = 8'hef;
        my_rom[3642] = 8'hef;
        my_rom[3643] = 8'hef;
        my_rom[3644] = 8'hf7;
        my_rom[3645] = 8'hf7;
        my_rom[3646] = 8'hef;
        my_rom[3647] = 8'hef;
        my_rom[3648] = 8'hf7;
        my_rom[3649] = 8'hef;
        my_rom[3650] = 8'hef;
        my_rom[3651] = 8'haf;
        my_rom[3652] = 8'had;
        my_rom[3653] = 8'ha5;
        my_rom[3654] = 8'ha5;
        my_rom[3655] = 8'ha5;
        my_rom[3656] = 8'ha5;
        my_rom[3657] = 8'ha5;
        my_rom[3658] = 8'ha5;
        my_rom[3659] = 8'haf;
        my_rom[3660] = 8'haf;
        my_rom[3661] = 8'had;
        my_rom[3662] = 8'ha5;
        my_rom[3663] = 8'h53;
        my_rom[3664] = 8'h49;
        my_rom[3665] = 8'h49;
        my_rom[3666] = 8'h49;
        my_rom[3667] = 8'h5b;
        my_rom[3668] = 8'h8;
        my_rom[3669] = 8'h8;
        my_rom[3670] = 8'h8;
        my_rom[3671] = 8'ha;
        my_rom[3672] = 8'h8;
        my_rom[3673] = 8'h8;
        my_rom[3674] = 8'had;
        my_rom[3675] = 8'h5b;
        my_rom[3676] = 8'h53;
        my_rom[3677] = 8'h53;
        my_rom[3678] = 8'h53;
        my_rom[3679] = 8'h53;
        my_rom[3680] = 8'h53;
        my_rom[3681] = 8'h49;
        my_rom[3682] = 8'h49;
        my_rom[3683] = 8'h53;
        my_rom[3684] = 8'ha5;
        my_rom[3685] = 8'hf7;
        my_rom[3686] = 8'hf7;
        my_rom[3687] = 8'hf7;
        my_rom[3688] = 8'hf7;
        my_rom[3689] = 8'hf7;
        my_rom[3690] = 8'ha5;
        my_rom[3691] = 8'h9d;
        my_rom[3692] = 8'h5b;
        my_rom[3693] = 8'h53;
        my_rom[3694] = 8'h53;
        my_rom[3695] = 8'h53;
        my_rom[3696] = 8'h4b;
        my_rom[3697] = 8'h53;
        my_rom[3698] = 8'h53;
        my_rom[3699] = 8'h53;
        my_rom[3700] = 8'h5b;
        my_rom[3701] = 8'h9d;
        my_rom[3702] = 8'ha5;
        my_rom[3703] = 8'hef;
        my_rom[3704] = 8'hef;
        my_rom[3705] = 8'hef;
        my_rom[3706] = 8'hef;
        my_rom[3707] = 8'hef;
        my_rom[3708] = 8'hef;
        my_rom[3709] = 8'had;
        my_rom[3710] = 8'ha5;
        my_rom[3711] = 8'h9d;
        my_rom[3712] = 8'h53;
        my_rom[3713] = 8'h4b;
        my_rom[3714] = 8'hb;
        my_rom[3715] = 8'hb;
        my_rom[3716] = 8'hb;
        my_rom[3717] = 8'hb;
        my_rom[3718] = 8'h53;
        my_rom[3719] = 8'h5b;
        my_rom[3720] = 8'ha5;
        my_rom[3721] = 8'had;
        my_rom[3722] = 8'had;
        my_rom[3723] = 8'h53;
        my_rom[3724] = 8'h49;
        my_rom[3725] = 8'h49;
        my_rom[3726] = 8'h51;
        my_rom[3727] = 8'h9b;
        my_rom[3728] = 8'h8;
        my_rom[3729] = 8'h8;
        my_rom[3730] = 8'h8;
        my_rom[3731] = 8'ha;
        my_rom[3732] = 8'h8;
        my_rom[3733] = 8'h8;
        my_rom[3734] = 8'hed;
        my_rom[3735] = 8'h5b;
        my_rom[3736] = 8'h53;
        my_rom[3737] = 8'h53;
        my_rom[3738] = 8'h53;
        my_rom[3739] = 8'h53;
        my_rom[3740] = 8'h53;
        my_rom[3741] = 8'h9;
        my_rom[3742] = 8'h49;
        my_rom[3743] = 8'h5b;
        my_rom[3744] = 8'had;
        my_rom[3745] = 8'hf7;
        my_rom[3746] = 8'hf7;
        my_rom[3747] = 8'hf7;
        my_rom[3748] = 8'had;
        my_rom[3749] = 8'ha5;
        my_rom[3750] = 8'ha5;
        my_rom[3751] = 8'ha5;
        my_rom[3752] = 8'h9d;
        my_rom[3753] = 8'h9d;
        my_rom[3754] = 8'h9b;
        my_rom[3755] = 8'h53;
        my_rom[3756] = 8'h53;
        my_rom[3757] = 8'h53;
        my_rom[3758] = 8'h53;
        my_rom[3759] = 8'h53;
        my_rom[3760] = 8'h53;
        my_rom[3761] = 8'h53;
        my_rom[3762] = 8'ha5;
        my_rom[3763] = 8'had;
        my_rom[3764] = 8'hed;
        my_rom[3765] = 8'hed;
        my_rom[3766] = 8'hed;
        my_rom[3767] = 8'hed;
        my_rom[3768] = 8'ha5;
        my_rom[3769] = 8'ha5;
        my_rom[3770] = 8'h9b;
        my_rom[3771] = 8'h53;
        my_rom[3772] = 8'h4b;
        my_rom[3773] = 8'h49;
        my_rom[3774] = 8'h9;
        my_rom[3775] = 8'h9;
        my_rom[3776] = 8'h49;
        my_rom[3777] = 8'h4b;
        my_rom[3778] = 8'h4b;
        my_rom[3779] = 8'h53;
        my_rom[3780] = 8'h53;
        my_rom[3781] = 8'h5b;
        my_rom[3782] = 8'ha5;
        my_rom[3783] = 8'h53;
        my_rom[3784] = 8'h9;
        my_rom[3785] = 8'h49;
        my_rom[3786] = 8'h53;
        my_rom[3787] = 8'ha3;
        my_rom[3788] = 8'h8;
        my_rom[3789] = 8'h8;
        my_rom[3790] = 8'h8;
        my_rom[3791] = 8'ha;
        my_rom[3792] = 8'h8;
        my_rom[3793] = 8'h8;
        my_rom[3794] = 8'h8;
        my_rom[3795] = 8'h5b;
        my_rom[3796] = 8'h53;
        my_rom[3797] = 8'h53;
        my_rom[3798] = 8'h53;
        my_rom[3799] = 8'h53;
        my_rom[3800] = 8'h53;
        my_rom[3801] = 8'h49;
        my_rom[3802] = 8'h49;
        my_rom[3803] = 8'h9b;
        my_rom[3804] = 8'hed;
        my_rom[3805] = 8'hf7;
        my_rom[3806] = 8'hf7;
        my_rom[3807] = 8'hed;
        my_rom[3808] = 8'ha5;
        my_rom[3809] = 8'had;
        my_rom[3810] = 8'had;
        my_rom[3811] = 8'had;
        my_rom[3812] = 8'had;
        my_rom[3813] = 8'ha5;
        my_rom[3814] = 8'ha5;
        my_rom[3815] = 8'ha5;
        my_rom[3816] = 8'h9b;
        my_rom[3817] = 8'h9b;
        my_rom[3818] = 8'h9b;
        my_rom[3819] = 8'h9b;
        my_rom[3820] = 8'h9b;
        my_rom[3821] = 8'h9b;
        my_rom[3822] = 8'h9b;
        my_rom[3823] = 8'ha5;
        my_rom[3824] = 8'hed;
        my_rom[3825] = 8'hed;
        my_rom[3826] = 8'ha5;
        my_rom[3827] = 8'ha5;
        my_rom[3828] = 8'ha5;
        my_rom[3829] = 8'h9b;
        my_rom[3830] = 8'h9b;
        my_rom[3831] = 8'h9b;
        my_rom[3832] = 8'h93;
        my_rom[3833] = 8'h53;
        my_rom[3834] = 8'h53;
        my_rom[3835] = 8'h9b;
        my_rom[3836] = 8'h9b;
        my_rom[3837] = 8'h9b;
        my_rom[3838] = 8'h9b;
        my_rom[3839] = 8'h5b;
        my_rom[3840] = 8'h5b;
        my_rom[3841] = 8'h5b;
        my_rom[3842] = 8'ha5;
        my_rom[3843] = 8'h53;
        my_rom[3844] = 8'h9;
        my_rom[3845] = 8'h49;
        my_rom[3846] = 8'h53;
        my_rom[3847] = 8'ha3;
        my_rom[3848] = 8'h8;
        my_rom[3849] = 8'h8;
        my_rom[3850] = 8'h8;
        my_rom[3851] = 8'ha;
        my_rom[3852] = 8'h8;
        my_rom[3853] = 8'h8;
        my_rom[3854] = 8'h8;
        my_rom[3855] = 8'ha3;
        my_rom[3856] = 8'h53;
        my_rom[3857] = 8'h53;
        my_rom[3858] = 8'h53;
        my_rom[3859] = 8'h53;
        my_rom[3860] = 8'h4b;
        my_rom[3861] = 8'h49;
        my_rom[3862] = 8'h53;
        my_rom[3863] = 8'ha5;
        my_rom[3864] = 8'hf7;
        my_rom[3865] = 8'hf7;
        my_rom[3866] = 8'hf7;
        my_rom[3867] = 8'had;
        my_rom[3868] = 8'had;
        my_rom[3869] = 8'hed;
        my_rom[3870] = 8'hed;
        my_rom[3871] = 8'hed;
        my_rom[3872] = 8'hed;
        my_rom[3873] = 8'ha5;
        my_rom[3874] = 8'ha5;
        my_rom[3875] = 8'ha5;
        my_rom[3876] = 8'h9b;
        my_rom[3877] = 8'h9b;
        my_rom[3878] = 8'h9b;
        my_rom[3879] = 8'h9b;
        my_rom[3880] = 8'h9b;
        my_rom[3881] = 8'h9b;
        my_rom[3882] = 8'ha3;
        my_rom[3883] = 8'ha5;
        my_rom[3884] = 8'hed;
        my_rom[3885] = 8'hed;
        my_rom[3886] = 8'ha5;
        my_rom[3887] = 8'ha5;
        my_rom[3888] = 8'ha3;
        my_rom[3889] = 8'h9b;
        my_rom[3890] = 8'h9b;
        my_rom[3891] = 8'h9b;
        my_rom[3892] = 8'h9b;
        my_rom[3893] = 8'h93;
        my_rom[3894] = 8'h9b;
        my_rom[3895] = 8'h9b;
        my_rom[3896] = 8'h9b;
        my_rom[3897] = 8'h9b;
        my_rom[3898] = 8'ha5;
        my_rom[3899] = 8'ha5;
        my_rom[3900] = 8'ha5;
        my_rom[3901] = 8'h9d;
        my_rom[3902] = 8'ha5;
        my_rom[3903] = 8'h53;
        my_rom[3904] = 8'h9;
        my_rom[3905] = 8'h49;
        my_rom[3906] = 8'h53;
        my_rom[3907] = 8'ha3;
        my_rom[3908] = 8'h8;
        my_rom[3909] = 8'h8;
        my_rom[3910] = 8'h8;
        my_rom[3911] = 8'ha;
        my_rom[3912] = 8'h8;
        my_rom[3913] = 8'hf5;
        my_rom[3914] = 8'hf5;
        my_rom[3915] = 8'hf7;
        my_rom[3916] = 8'hed;
        my_rom[3917] = 8'h53;
        my_rom[3918] = 8'h53;
        my_rom[3919] = 8'h53;
        my_rom[3920] = 8'h4b;
        my_rom[3921] = 8'h49;
        my_rom[3922] = 8'h53;
        my_rom[3923] = 8'ha5;
        my_rom[3924] = 8'hf7;
        my_rom[3925] = 8'hf7;
        my_rom[3926] = 8'hf7;
        my_rom[3927] = 8'hed;
        my_rom[3928] = 8'hed;
        my_rom[3929] = 8'hed;
        my_rom[3930] = 8'hed;
        my_rom[3931] = 8'ha5;
        my_rom[3932] = 8'h9b;
        my_rom[3933] = 8'h9d;
        my_rom[3934] = 8'ha5;
        my_rom[3935] = 8'h9d;
        my_rom[3936] = 8'h53;
        my_rom[3937] = 8'h53;
        my_rom[3938] = 8'h49;
        my_rom[3939] = 8'h93;
        my_rom[3940] = 8'h9b;
        my_rom[3941] = 8'h9b;
        my_rom[3942] = 8'ha5;
        my_rom[3943] = 8'ha5;
        my_rom[3944] = 8'hed;
        my_rom[3945] = 8'hed;
        my_rom[3946] = 8'hed;
        my_rom[3947] = 8'ha5;
        my_rom[3948] = 8'ha3;
        my_rom[3949] = 8'h9b;
        my_rom[3950] = 8'h9b;
        my_rom[3951] = 8'h93;
        my_rom[3952] = 8'h53;
        my_rom[3953] = 8'h49;
        my_rom[3954] = 8'h53;
        my_rom[3955] = 8'h53;
        my_rom[3956] = 8'h53;
        my_rom[3957] = 8'h53;
        my_rom[3958] = 8'h9b;
        my_rom[3959] = 8'h9b;
        my_rom[3960] = 8'ha5;
        my_rom[3961] = 8'ha5;
        my_rom[3962] = 8'ha5;
        my_rom[3963] = 8'h53;
        my_rom[3964] = 8'h9;
        my_rom[3965] = 8'h49;
        my_rom[3966] = 8'h53;
        my_rom[3967] = 8'ha3;
        my_rom[3968] = 8'ha3;
        my_rom[3969] = 8'h8;
        my_rom[3970] = 8'h8;
        my_rom[3971] = 8'ha;
        my_rom[3972] = 8'h8;
        my_rom[3973] = 8'hf5;
        my_rom[3974] = 8'hf7;
        my_rom[3975] = 8'hed;
        my_rom[3976] = 8'hed;
        my_rom[3977] = 8'h53;
        my_rom[3978] = 8'h53;
        my_rom[3979] = 8'h53;
        my_rom[3980] = 8'h4b;
        my_rom[3981] = 8'h49;
        my_rom[3982] = 8'h53;
        my_rom[3983] = 8'ha5;
        my_rom[3984] = 8'hf7;
        my_rom[3985] = 8'hf7;
        my_rom[3986] = 8'hf7;
        my_rom[3987] = 8'hf7;
        my_rom[3988] = 8'hed;
        my_rom[3989] = 8'hed;
        my_rom[3990] = 8'ha5;
        my_rom[3991] = 8'h9b;
        my_rom[3992] = 8'ha5;
        my_rom[3993] = 8'ha5;
        my_rom[3994] = 8'h5b;
        my_rom[3995] = 8'h53;
        my_rom[3996] = 8'h4b;
        my_rom[3997] = 8'h4b;
        my_rom[3998] = 8'h53;
        my_rom[3999] = 8'h53;
        my_rom[4000] = 8'h53;
        my_rom[4001] = 8'h9b;
        my_rom[4002] = 8'ha5;
        my_rom[4003] = 8'hed;
        my_rom[4004] = 8'hf7;
        my_rom[4005] = 8'hf7;
        my_rom[4006] = 8'hef;
        my_rom[4007] = 8'had;
        my_rom[4008] = 8'ha3;
        my_rom[4009] = 8'h9b;
        my_rom[4010] = 8'h93;
        my_rom[4011] = 8'h49;
        my_rom[4012] = 8'h49;
        my_rom[4013] = 8'h53;
        my_rom[4014] = 8'h53;
        my_rom[4015] = 8'h53;
        my_rom[4016] = 8'h5b;
        my_rom[4017] = 8'h9d;
        my_rom[4018] = 8'h9b;
        my_rom[4019] = 8'h93;
        my_rom[4020] = 8'ha3;
        my_rom[4021] = 8'ha5;
        my_rom[4022] = 8'had;
        my_rom[4023] = 8'h53;
        my_rom[4024] = 8'h9;
        my_rom[4025] = 8'h49;
        my_rom[4026] = 8'h9b;
        my_rom[4027] = 8'ha5;
        my_rom[4028] = 8'had;
        my_rom[4029] = 8'had;
        my_rom[4030] = 8'h8;
        my_rom[4031] = 8'ha;
        my_rom[4032] = 8'hf5;
        my_rom[4033] = 8'hf7;
        my_rom[4034] = 8'he5;
        my_rom[4035] = 8'h93;
        my_rom[4036] = 8'h9b;
        my_rom[4037] = 8'h53;
        my_rom[4038] = 8'h53;
        my_rom[4039] = 8'h53;
        my_rom[4040] = 8'h4b;
        my_rom[4041] = 8'h9;
        my_rom[4042] = 8'h53;
        my_rom[4043] = 8'had;
        my_rom[4044] = 8'hf7;
        my_rom[4045] = 8'hf7;
        my_rom[4046] = 8'hf7;
        my_rom[4047] = 8'hf7;
        my_rom[4048] = 8'hed;
        my_rom[4049] = 8'he5;
        my_rom[4050] = 8'h9b;
        my_rom[4051] = 8'ha5;
        my_rom[4052] = 8'h5b;
        my_rom[4053] = 8'h49;
        my_rom[4054] = 8'h9;
        my_rom[4055] = 8'h1;
        my_rom[4056] = 8'h49;
        my_rom[4057] = 8'h5b;
        my_rom[4058] = 8'h53;
        my_rom[4059] = 8'h4b;
        my_rom[4060] = 8'h53;
        my_rom[4061] = 8'h9b;
        my_rom[4062] = 8'ha5;
        my_rom[4063] = 8'hed;
        my_rom[4064] = 8'hf7;
        my_rom[4065] = 8'hf7;
        my_rom[4066] = 8'hf7;
        my_rom[4067] = 8'had;
        my_rom[4068] = 8'ha5;
        my_rom[4069] = 8'h9b;
        my_rom[4070] = 8'h53;
        my_rom[4071] = 8'h49;
        my_rom[4072] = 8'h49;
        my_rom[4073] = 8'h9;
        my_rom[4074] = 8'h9;
        my_rom[4075] = 8'h9;
        my_rom[4076] = 8'h9;
        my_rom[4077] = 8'h53;
        my_rom[4078] = 8'h9d;
        my_rom[4079] = 8'h9b;
        my_rom[4080] = 8'h9b;
        my_rom[4081] = 8'ha5;
        my_rom[4082] = 8'had;
        my_rom[4083] = 8'h5b;
        my_rom[4084] = 8'h9;
        my_rom[4085] = 8'h53;
        my_rom[4086] = 8'ha5;
        my_rom[4087] = 8'hef;
        my_rom[4088] = 8'hed;
        my_rom[4089] = 8'had;
        my_rom[4090] = 8'h8;
        my_rom[4091] = 8'ha;
        my_rom[4092] = 8'hf5;
        my_rom[4093] = 8'hf5;
        my_rom[4094] = 8'hdb;
        my_rom[4095] = 8'hdb;
        my_rom[4096] = 8'hed;
        my_rom[4097] = 8'ha5;
        my_rom[4098] = 8'h9b;
        my_rom[4099] = 8'h5b;
        my_rom[4100] = 8'h53;
        my_rom[4101] = 8'h9;
        my_rom[4102] = 8'h49;
        my_rom[4103] = 8'had;
        my_rom[4104] = 8'hf7;
        my_rom[4105] = 8'hf7;
        my_rom[4106] = 8'hf7;
        my_rom[4107] = 8'hf7;
        my_rom[4108] = 8'hed;
        my_rom[4109] = 8'ha5;
        my_rom[4110] = 8'h9b;
        my_rom[4111] = 8'h53;
        my_rom[4112] = 8'h53;
        my_rom[4113] = 8'h5b;
        my_rom[4114] = 8'h53;
        my_rom[4115] = 8'h4b;
        my_rom[4116] = 8'h53;
        my_rom[4117] = 8'h9d;
        my_rom[4118] = 8'h9d;
        my_rom[4119] = 8'h53;
        my_rom[4120] = 8'h53;
        my_rom[4121] = 8'ha5;
        my_rom[4122] = 8'had;
        my_rom[4123] = 8'hf7;
        my_rom[4124] = 8'hf7;
        my_rom[4125] = 8'hf7;
        my_rom[4126] = 8'hf7;
        my_rom[4127] = 8'hef;
        my_rom[4128] = 8'ha5;
        my_rom[4129] = 8'h9b;
        my_rom[4130] = 8'h53;
        my_rom[4131] = 8'h53;
        my_rom[4132] = 8'h53;
        my_rom[4133] = 8'h49;
        my_rom[4134] = 8'h9;
        my_rom[4135] = 8'h49;
        my_rom[4136] = 8'h53;
        my_rom[4137] = 8'h53;
        my_rom[4138] = 8'h49;
        my_rom[4139] = 8'h5b;
        my_rom[4140] = 8'h9b;
        my_rom[4141] = 8'ha5;
        my_rom[4142] = 8'hed;
        my_rom[4143] = 8'h5b;
        my_rom[4144] = 8'h9;
        my_rom[4145] = 8'h53;
        my_rom[4146] = 8'h9b;
        my_rom[4147] = 8'h9b;
        my_rom[4148] = 8'he5;
        my_rom[4149] = 8'hf5;
        my_rom[4150] = 8'hf5;
        my_rom[4151] = 8'ha;
        my_rom[4152] = 8'hf5;
        my_rom[4153] = 8'hed;
        my_rom[4154] = 8'hdb;
        my_rom[4155] = 8'hed;
        my_rom[4156] = 8'hf7;
        my_rom[4157] = 8'hf7;
        my_rom[4158] = 8'ha5;
        my_rom[4159] = 8'h9b;
        my_rom[4160] = 8'h53;
        my_rom[4161] = 8'h9;
        my_rom[4162] = 8'h4b;
        my_rom[4163] = 8'had;
        my_rom[4164] = 8'hf7;
        my_rom[4165] = 8'hf7;
        my_rom[4166] = 8'hf7;
        my_rom[4167] = 8'hf7;
        my_rom[4168] = 8'hed;
        my_rom[4169] = 8'hed;
        my_rom[4170] = 8'hed;
        my_rom[4171] = 8'hed;
        my_rom[4172] = 8'ha5;
        my_rom[4173] = 8'ha5;
        my_rom[4174] = 8'h9d;
        my_rom[4175] = 8'h9d;
        my_rom[4176] = 8'h9d;
        my_rom[4177] = 8'h9d;
        my_rom[4178] = 8'h9d;
        my_rom[4179] = 8'h9d;
        my_rom[4180] = 8'ha5;
        my_rom[4181] = 8'ha5;
        my_rom[4182] = 8'hf7;
        my_rom[4183] = 8'hf7;
        my_rom[4184] = 8'hf7;
        my_rom[4185] = 8'hf7;
        my_rom[4186] = 8'hf7;
        my_rom[4187] = 8'hef;
        my_rom[4188] = 8'ha5;
        my_rom[4189] = 8'h9d;
        my_rom[4190] = 8'h9d;
        my_rom[4191] = 8'h9b;
        my_rom[4192] = 8'h9b;
        my_rom[4193] = 8'h5b;
        my_rom[4194] = 8'h53;
        my_rom[4195] = 8'h53;
        my_rom[4196] = 8'h53;
        my_rom[4197] = 8'h53;
        my_rom[4198] = 8'h53;
        my_rom[4199] = 8'h9b;
        my_rom[4200] = 8'h9d;
        my_rom[4201] = 8'ha5;
        my_rom[4202] = 8'hed;
        my_rom[4203] = 8'ha5;
        my_rom[4204] = 8'h49;
        my_rom[4205] = 8'h9b;
        my_rom[4206] = 8'h9b;
        my_rom[4207] = 8'h9b;
        my_rom[4208] = 8'h93;
        my_rom[4209] = 8'hed;
        my_rom[4210] = 8'hf5;
        my_rom[4211] = 8'ha;
        my_rom[4212] = 8'hf7;
        my_rom[4213] = 8'he5;
        my_rom[4214] = 8'hdb;
        my_rom[4215] = 8'hed;
        my_rom[4216] = 8'hf7;
        my_rom[4217] = 8'hf7;
        my_rom[4218] = 8'hf7;
        my_rom[4219] = 8'h9b;
        my_rom[4220] = 8'h5b;
        my_rom[4221] = 8'h53;
        my_rom[4222] = 8'h53;
        my_rom[4223] = 8'hed;
        my_rom[4224] = 8'hf7;
        my_rom[4225] = 8'hf7;
        my_rom[4226] = 8'hf7;
        my_rom[4227] = 8'hf7;
        my_rom[4228] = 8'hf7;
        my_rom[4229] = 8'hf7;
        my_rom[4230] = 8'hf7;
        my_rom[4231] = 8'hed;
        my_rom[4232] = 8'hed;
        my_rom[4233] = 8'ha5;
        my_rom[4234] = 8'ha5;
        my_rom[4235] = 8'ha5;
        my_rom[4236] = 8'h9d;
        my_rom[4237] = 8'h9d;
        my_rom[4238] = 8'ha5;
        my_rom[4239] = 8'ha5;
        my_rom[4240] = 8'had;
        my_rom[4241] = 8'hf7;
        my_rom[4242] = 8'hf7;
        my_rom[4243] = 8'hf7;
        my_rom[4244] = 8'hf7;
        my_rom[4245] = 8'hff;
        my_rom[4246] = 8'hf7;
        my_rom[4247] = 8'hef;
        my_rom[4248] = 8'had;
        my_rom[4249] = 8'ha5;
        my_rom[4250] = 8'ha5;
        my_rom[4251] = 8'h9d;
        my_rom[4252] = 8'h9d;
        my_rom[4253] = 8'h9b;
        my_rom[4254] = 8'h9b;
        my_rom[4255] = 8'h9b;
        my_rom[4256] = 8'h9b;
        my_rom[4257] = 8'h9b;
        my_rom[4258] = 8'ha5;
        my_rom[4259] = 8'ha5;
        my_rom[4260] = 8'had;
        my_rom[4261] = 8'had;
        my_rom[4262] = 8'hef;
        my_rom[4263] = 8'ha5;
        my_rom[4264] = 8'h53;
        my_rom[4265] = 8'h9b;
        my_rom[4266] = 8'ha5;
        my_rom[4267] = 8'h9b;
        my_rom[4268] = 8'h93;
        my_rom[4269] = 8'hed;
        my_rom[4270] = 8'hf5;
        my_rom[4271] = 8'ha;
        my_rom[4272] = 8'hf7;
        my_rom[4273] = 8'he5;
        my_rom[4274] = 8'hdb;
        my_rom[4275] = 8'hef;
        my_rom[4276] = 8'hf7;
        my_rom[4277] = 8'hf7;
        my_rom[4278] = 8'hed;
        my_rom[4279] = 8'h9b;
        my_rom[4280] = 8'h9b;
        my_rom[4281] = 8'h53;
        my_rom[4282] = 8'h53;
        my_rom[4283] = 8'hed;
        my_rom[4284] = 8'hf7;
        my_rom[4285] = 8'hf7;
        my_rom[4286] = 8'hf7;
        my_rom[4287] = 8'hf7;
        my_rom[4288] = 8'hf7;
        my_rom[4289] = 8'hf7;
        my_rom[4290] = 8'hf7;
        my_rom[4291] = 8'hf7;
        my_rom[4292] = 8'hef;
        my_rom[4293] = 8'hed;
        my_rom[4294] = 8'hed;
        my_rom[4295] = 8'ha5;
        my_rom[4296] = 8'ha5;
        my_rom[4297] = 8'ha5;
        my_rom[4298] = 8'haf;
        my_rom[4299] = 8'haf;
        my_rom[4300] = 8'hf7;
        my_rom[4301] = 8'hf7;
        my_rom[4302] = 8'hf7;
        my_rom[4303] = 8'hf7;
        my_rom[4304] = 8'hf7;
        my_rom[4305] = 8'hff;
        my_rom[4306] = 8'hf7;
        my_rom[4307] = 8'hf7;
        my_rom[4308] = 8'hef;
        my_rom[4309] = 8'ha5;
        my_rom[4310] = 8'ha5;
        my_rom[4311] = 8'ha5;
        my_rom[4312] = 8'ha5;
        my_rom[4313] = 8'h9d;
        my_rom[4314] = 8'h9d;
        my_rom[4315] = 8'h9d;
        my_rom[4316] = 8'h9b;
        my_rom[4317] = 8'ha5;
        my_rom[4318] = 8'ha5;
        my_rom[4319] = 8'had;
        my_rom[4320] = 8'haf;
        my_rom[4321] = 8'hef;
        my_rom[4322] = 8'hef;
        my_rom[4323] = 8'ha5;
        my_rom[4324] = 8'h53;
        my_rom[4325] = 8'h9b;
        my_rom[4326] = 8'he5;
        my_rom[4327] = 8'hdd;
        my_rom[4328] = 8'h93;
        my_rom[4329] = 8'hed;
        my_rom[4330] = 8'hf5;
        my_rom[4331] = 8'ha;
        my_rom[4332] = 8'hf5;
        my_rom[4333] = 8'he5;
        my_rom[4334] = 8'he5;
        my_rom[4335] = 8'hf7;
        my_rom[4336] = 8'hf7;
        my_rom[4337] = 8'hed;
        my_rom[4338] = 8'h9b;
        my_rom[4339] = 8'h93;
        my_rom[4340] = 8'hed;
        my_rom[4341] = 8'h53;
        my_rom[4342] = 8'h53;
        my_rom[4343] = 8'hed;
        my_rom[4344] = 8'hf7;
        my_rom[4345] = 8'hf7;
        my_rom[4346] = 8'hf7;
        my_rom[4347] = 8'hf7;
        my_rom[4348] = 8'hf7;
        my_rom[4349] = 8'hf7;
        my_rom[4350] = 8'hf7;
        my_rom[4351] = 8'hf7;
        my_rom[4352] = 8'hf7;
        my_rom[4353] = 8'hf7;
        my_rom[4354] = 8'hef;
        my_rom[4355] = 8'hef;
        my_rom[4356] = 8'hef;
        my_rom[4357] = 8'hef;
        my_rom[4358] = 8'hf7;
        my_rom[4359] = 8'hf7;
        my_rom[4360] = 8'hf7;
        my_rom[4361] = 8'hf7;
        my_rom[4362] = 8'hf7;
        my_rom[4363] = 8'hf7;
        my_rom[4364] = 8'hf7;
        my_rom[4365] = 8'hff;
        my_rom[4366] = 8'hf7;
        my_rom[4367] = 8'hf7;
        my_rom[4368] = 8'hef;
        my_rom[4369] = 8'had;
        my_rom[4370] = 8'had;
        my_rom[4371] = 8'had;
        my_rom[4372] = 8'ha5;
        my_rom[4373] = 8'ha5;
        my_rom[4374] = 8'ha5;
        my_rom[4375] = 8'ha5;
        my_rom[4376] = 8'ha5;
        my_rom[4377] = 8'ha5;
        my_rom[4378] = 8'had;
        my_rom[4379] = 8'haf;
        my_rom[4380] = 8'hef;
        my_rom[4381] = 8'hef;
        my_rom[4382] = 8'hf7;
        my_rom[4383] = 8'had;
        my_rom[4384] = 8'h53;
        my_rom[4385] = 8'ha5;
        my_rom[4386] = 8'hed;
        my_rom[4387] = 8'he5;
        my_rom[4388] = 8'h9b;
        my_rom[4389] = 8'hed;
        my_rom[4390] = 8'h8;
        my_rom[4391] = 8'ha;
        my_rom[4392] = 8'hf7;
        my_rom[4393] = 8'hed;
        my_rom[4394] = 8'he5;
        my_rom[4395] = 8'hf7;
        my_rom[4396] = 8'hf7;
        my_rom[4397] = 8'he5;
        my_rom[4398] = 8'h9b;
        my_rom[4399] = 8'he5;
        my_rom[4400] = 8'hf7;
        my_rom[4401] = 8'ha5;
        my_rom[4402] = 8'h53;
        my_rom[4403] = 8'hf5;
        my_rom[4404] = 8'hf7;
        my_rom[4405] = 8'hf7;
        my_rom[4406] = 8'hf7;
        my_rom[4407] = 8'hf7;
        my_rom[4408] = 8'hf7;
        my_rom[4409] = 8'hf7;
        my_rom[4410] = 8'hf7;
        my_rom[4411] = 8'hf7;
        my_rom[4412] = 8'hf7;
        my_rom[4413] = 8'hf7;
        my_rom[4414] = 8'hf7;
        my_rom[4415] = 8'hf7;
        my_rom[4416] = 8'hf7;
        my_rom[4417] = 8'hf7;
        my_rom[4418] = 8'hf7;
        my_rom[4419] = 8'hf7;
        my_rom[4420] = 8'hf7;
        my_rom[4421] = 8'hf7;
        my_rom[4422] = 8'hf7;
        my_rom[4423] = 8'hf7;
        my_rom[4424] = 8'hf7;
        my_rom[4425] = 8'hf7;
        my_rom[4426] = 8'hf7;
        my_rom[4427] = 8'hf7;
        my_rom[4428] = 8'hef;
        my_rom[4429] = 8'hef;
        my_rom[4430] = 8'had;
        my_rom[4431] = 8'had;
        my_rom[4432] = 8'haf;
        my_rom[4433] = 8'haf;
        my_rom[4434] = 8'had;
        my_rom[4435] = 8'had;
        my_rom[4436] = 8'had;
        my_rom[4437] = 8'haf;
        my_rom[4438] = 8'haf;
        my_rom[4439] = 8'hef;
        my_rom[4440] = 8'hef;
        my_rom[4441] = 8'hf7;
        my_rom[4442] = 8'hf7;
        my_rom[4443] = 8'had;
        my_rom[4444] = 8'h93;
        my_rom[4445] = 8'h9b;
        my_rom[4446] = 8'hed;
        my_rom[4447] = 8'he5;
        my_rom[4448] = 8'h9b;
        my_rom[4449] = 8'hed;
        my_rom[4450] = 8'h8;
        my_rom[4451] = 8'ha;
        my_rom[4452] = 8'hf5;
        my_rom[4453] = 8'hf7;
        my_rom[4454] = 8'hed;
        my_rom[4455] = 8'hf7;
        my_rom[4456] = 8'hed;
        my_rom[4457] = 8'he3;
        my_rom[4458] = 8'h9b;
        my_rom[4459] = 8'hed;
        my_rom[4460] = 8'hf7;
        my_rom[4461] = 8'ha5;
        my_rom[4462] = 8'h53;
        my_rom[4463] = 8'hf7;
        my_rom[4464] = 8'hf7;
        my_rom[4465] = 8'hf7;
        my_rom[4466] = 8'hf7;
        my_rom[4467] = 8'hf7;
        my_rom[4468] = 8'hf7;
        my_rom[4469] = 8'hf7;
        my_rom[4470] = 8'hf7;
        my_rom[4471] = 8'hf7;
        my_rom[4472] = 8'hf7;
        my_rom[4473] = 8'hf7;
        my_rom[4474] = 8'hf7;
        my_rom[4475] = 8'hf7;
        my_rom[4476] = 8'hf7;
        my_rom[4477] = 8'hf7;
        my_rom[4478] = 8'hf7;
        my_rom[4479] = 8'hf7;
        my_rom[4480] = 8'hf7;
        my_rom[4481] = 8'hf7;
        my_rom[4482] = 8'hf7;
        my_rom[4483] = 8'hf7;
        my_rom[4484] = 8'hf7;
        my_rom[4485] = 8'hf7;
        my_rom[4486] = 8'hf7;
        my_rom[4487] = 8'hf7;
        my_rom[4488] = 8'hf7;
        my_rom[4489] = 8'hef;
        my_rom[4490] = 8'haf;
        my_rom[4491] = 8'haf;
        my_rom[4492] = 8'haf;
        my_rom[4493] = 8'haf;
        my_rom[4494] = 8'haf;
        my_rom[4495] = 8'haf;
        my_rom[4496] = 8'haf;
        my_rom[4497] = 8'haf;
        my_rom[4498] = 8'hef;
        my_rom[4499] = 8'hef;
        my_rom[4500] = 8'hf7;
        my_rom[4501] = 8'hf7;
        my_rom[4502] = 8'hef;
        my_rom[4503] = 8'had;
        my_rom[4504] = 8'h93;
        my_rom[4505] = 8'h9b;
        my_rom[4506] = 8'ha5;
        my_rom[4507] = 8'he5;
        my_rom[4508] = 8'he5;
        my_rom[4509] = 8'hed;
        my_rom[4510] = 8'h8;
        my_rom[4511] = 8'ha;
        my_rom[4512] = 8'h8;
        my_rom[4513] = 8'hf7;
        my_rom[4514] = 8'hf7;
        my_rom[4515] = 8'hf7;
        my_rom[4516] = 8'hed;
        my_rom[4517] = 8'he5;
        my_rom[4518] = 8'he5;
        my_rom[4519] = 8'hed;
        my_rom[4520] = 8'hed;
        my_rom[4521] = 8'hed;
        my_rom[4522] = 8'h9b;
        my_rom[4523] = 8'hf5;
        my_rom[4524] = 8'hf7;
        my_rom[4525] = 8'hf7;
        my_rom[4526] = 8'hf7;
        my_rom[4527] = 8'hf7;
        my_rom[4528] = 8'hf7;
        my_rom[4529] = 8'hf7;
        my_rom[4530] = 8'hf7;
        my_rom[4531] = 8'hf7;
        my_rom[4532] = 8'hf7;
        my_rom[4533] = 8'hf7;
        my_rom[4534] = 8'hf7;
        my_rom[4535] = 8'hf7;
        my_rom[4536] = 8'hf7;
        my_rom[4537] = 8'hf7;
        my_rom[4538] = 8'hf7;
        my_rom[4539] = 8'hf7;
        my_rom[4540] = 8'hf7;
        my_rom[4541] = 8'hf7;
        my_rom[4542] = 8'hf7;
        my_rom[4543] = 8'hf7;
        my_rom[4544] = 8'hf7;
        my_rom[4545] = 8'hf7;
        my_rom[4546] = 8'hf7;
        my_rom[4547] = 8'hf7;
        my_rom[4548] = 8'hf7;
        my_rom[4549] = 8'hef;
        my_rom[4550] = 8'haf;
        my_rom[4551] = 8'haf;
        my_rom[4552] = 8'hef;
        my_rom[4553] = 8'hef;
        my_rom[4554] = 8'hef;
        my_rom[4555] = 8'hef;
        my_rom[4556] = 8'hef;
        my_rom[4557] = 8'hef;
        my_rom[4558] = 8'hef;
        my_rom[4559] = 8'hf7;
        my_rom[4560] = 8'hf7;
        my_rom[4561] = 8'hef;
        my_rom[4562] = 8'hef;
        my_rom[4563] = 8'hef;
        my_rom[4564] = 8'h93;
        my_rom[4565] = 8'h9b;
        my_rom[4566] = 8'ha5;
        my_rom[4567] = 8'hed;
        my_rom[4568] = 8'hed;
        my_rom[4569] = 8'hf5;
        my_rom[4570] = 8'h8;
        my_rom[4571] = 8'ha;
        my_rom[4572] = 8'h8;
        my_rom[4573] = 8'hf5;
        my_rom[4574] = 8'hf7;
        my_rom[4575] = 8'hef;
        my_rom[4576] = 8'hef;
        my_rom[4577] = 8'he5;
        my_rom[4578] = 8'he5;
        my_rom[4579] = 8'he5;
        my_rom[4580] = 8'hed;
        my_rom[4581] = 8'hf7;
        my_rom[4582] = 8'hed;
        my_rom[4583] = 8'hf7;
        my_rom[4584] = 8'hf7;
        my_rom[4585] = 8'hf7;
        my_rom[4586] = 8'hf7;
        my_rom[4587] = 8'hf7;
        my_rom[4588] = 8'hf7;
        my_rom[4589] = 8'hf7;
        my_rom[4590] = 8'hf7;
        my_rom[4591] = 8'hf7;
        my_rom[4592] = 8'hf7;
        my_rom[4593] = 8'hf7;
        my_rom[4594] = 8'hf7;
        my_rom[4595] = 8'hf7;
        my_rom[4596] = 8'hf7;
        my_rom[4597] = 8'hf7;
        my_rom[4598] = 8'hf7;
        my_rom[4599] = 8'hf7;
        my_rom[4600] = 8'hf7;
        my_rom[4601] = 8'hf7;
        my_rom[4602] = 8'hf7;
        my_rom[4603] = 8'hf7;
        my_rom[4604] = 8'hf7;
        my_rom[4605] = 8'hf7;
        my_rom[4606] = 8'hf7;
        my_rom[4607] = 8'hf7;
        my_rom[4608] = 8'hef;
        my_rom[4609] = 8'hef;
        my_rom[4610] = 8'hef;
        my_rom[4611] = 8'had;
        my_rom[4612] = 8'hef;
        my_rom[4613] = 8'haf;
        my_rom[4614] = 8'hef;
        my_rom[4615] = 8'hef;
        my_rom[4616] = 8'hef;
        my_rom[4617] = 8'hef;
        my_rom[4618] = 8'hef;
        my_rom[4619] = 8'hef;
        my_rom[4620] = 8'hef;
        my_rom[4621] = 8'hef;
        my_rom[4622] = 8'hef;
        my_rom[4623] = 8'hed;
        my_rom[4624] = 8'h93;
        my_rom[4625] = 8'h9b;
        my_rom[4626] = 8'ha5;
        my_rom[4627] = 8'he5;
        my_rom[4628] = 8'hed;
        my_rom[4629] = 8'h8;
        my_rom[4630] = 8'h8;
        my_rom[4631] = 8'ha;
        my_rom[4632] = 8'h8;
        my_rom[4633] = 8'hf5;
        my_rom[4634] = 8'hf7;
        my_rom[4635] = 8'hf7;
        my_rom[4636] = 8'hed;
        my_rom[4637] = 8'hed;
        my_rom[4638] = 8'he5;
        my_rom[4639] = 8'hed;
        my_rom[4640] = 8'hef;
        my_rom[4641] = 8'hf7;
        my_rom[4642] = 8'hf7;
        my_rom[4643] = 8'hf7;
        my_rom[4644] = 8'hf7;
        my_rom[4645] = 8'hf7;
        my_rom[4646] = 8'hf7;
        my_rom[4647] = 8'hf7;
        my_rom[4648] = 8'hf7;
        my_rom[4649] = 8'hf7;
        my_rom[4650] = 8'hf7;
        my_rom[4651] = 8'hf7;
        my_rom[4652] = 8'hf7;
        my_rom[4653] = 8'hf7;
        my_rom[4654] = 8'hf7;
        my_rom[4655] = 8'hf7;
        my_rom[4656] = 8'hf7;
        my_rom[4657] = 8'hf7;
        my_rom[4658] = 8'hef;
        my_rom[4659] = 8'hef;
        my_rom[4660] = 8'hf7;
        my_rom[4661] = 8'hf7;
        my_rom[4662] = 8'hf7;
        my_rom[4663] = 8'hf7;
        my_rom[4664] = 8'hf7;
        my_rom[4665] = 8'hf7;
        my_rom[4666] = 8'hf7;
        my_rom[4667] = 8'hef;
        my_rom[4668] = 8'hef;
        my_rom[4669] = 8'hef;
        my_rom[4670] = 8'hef;
        my_rom[4671] = 8'had;
        my_rom[4672] = 8'haf;
        my_rom[4673] = 8'hef;
        my_rom[4674] = 8'hef;
        my_rom[4675] = 8'hef;
        my_rom[4676] = 8'hef;
        my_rom[4677] = 8'hef;
        my_rom[4678] = 8'hef;
        my_rom[4679] = 8'hef;
        my_rom[4680] = 8'hef;
        my_rom[4681] = 8'hef;
        my_rom[4682] = 8'hef;
        my_rom[4683] = 8'hed;
        my_rom[4684] = 8'h93;
        my_rom[4685] = 8'h9d;
        my_rom[4686] = 8'ha5;
        my_rom[4687] = 8'he5;
        my_rom[4688] = 8'hed;
        my_rom[4689] = 8'h8;
        my_rom[4690] = 8'h8;
        my_rom[4691] = 8'ha;
        my_rom[4692] = 8'h8;
        my_rom[4693] = 8'hf5;
        my_rom[4694] = 8'hf5;
        my_rom[4695] = 8'hf7;
        my_rom[4696] = 8'hed;
        my_rom[4697] = 8'hed;
        my_rom[4698] = 8'hf7;
        my_rom[4699] = 8'hf7;
        my_rom[4700] = 8'hf7;
        my_rom[4701] = 8'hf7;
        my_rom[4702] = 8'hf7;
        my_rom[4703] = 8'hf7;
        my_rom[4704] = 8'hf7;
        my_rom[4705] = 8'hf7;
        my_rom[4706] = 8'hf7;
        my_rom[4707] = 8'hf7;
        my_rom[4708] = 8'hf7;
        my_rom[4709] = 8'hf7;
        my_rom[4710] = 8'hf7;
        my_rom[4711] = 8'hf7;
        my_rom[4712] = 8'hf7;
        my_rom[4713] = 8'hf7;
        my_rom[4714] = 8'hf7;
        my_rom[4715] = 8'hf7;
        my_rom[4716] = 8'hf7;
        my_rom[4717] = 8'hef;
        my_rom[4718] = 8'hed;
        my_rom[4719] = 8'hed;
        my_rom[4720] = 8'hf7;
        my_rom[4721] = 8'hf7;
        my_rom[4722] = 8'hf7;
        my_rom[4723] = 8'hed;
        my_rom[4724] = 8'hed;
        my_rom[4725] = 8'hed;
        my_rom[4726] = 8'he5;
        my_rom[4727] = 8'ha5;
        my_rom[4728] = 8'ha5;
        my_rom[4729] = 8'he5;
        my_rom[4730] = 8'he5;
        my_rom[4731] = 8'hef;
        my_rom[4732] = 8'ha5;
        my_rom[4733] = 8'haf;
        my_rom[4734] = 8'hef;
        my_rom[4735] = 8'hef;
        my_rom[4736] = 8'hef;
        my_rom[4737] = 8'hef;
        my_rom[4738] = 8'hef;
        my_rom[4739] = 8'hef;
        my_rom[4740] = 8'hef;
        my_rom[4741] = 8'hef;
        my_rom[4742] = 8'hed;
        my_rom[4743] = 8'had;
        my_rom[4744] = 8'h9d;
        my_rom[4745] = 8'ha5;
        my_rom[4746] = 8'h9d;
        my_rom[4747] = 8'hed;
        my_rom[4748] = 8'hf5;
        my_rom[4749] = 8'h8;
        my_rom[4750] = 8'h8;
        my_rom[4751] = 8'ha;
        my_rom[4752] = 8'h8;
        my_rom[4753] = 8'h8;
        my_rom[4754] = 8'hf5;
        my_rom[4755] = 8'hf7;
        my_rom[4756] = 8'hf7;
        my_rom[4757] = 8'hf7;
        my_rom[4758] = 8'hf7;
        my_rom[4759] = 8'hf7;
        my_rom[4760] = 8'hf7;
        my_rom[4761] = 8'hf7;
        my_rom[4762] = 8'hf7;
        my_rom[4763] = 8'hf7;
        my_rom[4764] = 8'hf7;
        my_rom[4765] = 8'hf7;
        my_rom[4766] = 8'hf7;
        my_rom[4767] = 8'hf7;
        my_rom[4768] = 8'hf7;
        my_rom[4769] = 8'hf7;
        my_rom[4770] = 8'hf7;
        my_rom[4771] = 8'hf7;
        my_rom[4772] = 8'hf7;
        my_rom[4773] = 8'hf7;
        my_rom[4774] = 8'hf7;
        my_rom[4775] = 8'hf7;
        my_rom[4776] = 8'hef;
        my_rom[4777] = 8'hed;
        my_rom[4778] = 8'hed;
        my_rom[4779] = 8'hed;
        my_rom[4780] = 8'hef;
        my_rom[4781] = 8'hef;
        my_rom[4782] = 8'he5;
        my_rom[4783] = 8'h9b;
        my_rom[4784] = 8'h9b;
        my_rom[4785] = 8'ha5;
        my_rom[4786] = 8'h9b;
        my_rom[4787] = 8'h9b;
        my_rom[4788] = 8'h9b;
        my_rom[4789] = 8'h9b;
        my_rom[4790] = 8'h9b;
        my_rom[4791] = 8'he5;
        my_rom[4792] = 8'ha5;
        my_rom[4793] = 8'had;
        my_rom[4794] = 8'hef;
        my_rom[4795] = 8'hef;
        my_rom[4796] = 8'hef;
        my_rom[4797] = 8'hef;
        my_rom[4798] = 8'hef;
        my_rom[4799] = 8'hef;
        my_rom[4800] = 8'hef;
        my_rom[4801] = 8'hef;
        my_rom[4802] = 8'hed;
        my_rom[4803] = 8'hef;
        my_rom[4804] = 8'had;
        my_rom[4805] = 8'h9d;
        my_rom[4806] = 8'ha5;
        my_rom[4807] = 8'hed;
        my_rom[4808] = 8'hf5;
        my_rom[4809] = 8'h8;
        my_rom[4810] = 8'h8;
        my_rom[4811] = 8'ha;
        my_rom[4812] = 8'h8;
        my_rom[4813] = 8'h8;
        my_rom[4814] = 8'hf5;
        my_rom[4815] = 8'hf7;
        my_rom[4816] = 8'hf7;
        my_rom[4817] = 8'hf7;
        my_rom[4818] = 8'hff;
        my_rom[4819] = 8'hf7;
        my_rom[4820] = 8'hf7;
        my_rom[4821] = 8'hf7;
        my_rom[4822] = 8'hf7;
        my_rom[4823] = 8'hf7;
        my_rom[4824] = 8'hf7;
        my_rom[4825] = 8'hf7;
        my_rom[4826] = 8'hf7;
        my_rom[4827] = 8'hf7;
        my_rom[4828] = 8'hf7;
        my_rom[4829] = 8'hf7;
        my_rom[4830] = 8'hf7;
        my_rom[4831] = 8'hf7;
        my_rom[4832] = 8'hf7;
        my_rom[4833] = 8'hf7;
        my_rom[4834] = 8'hf7;
        my_rom[4835] = 8'hef;
        my_rom[4836] = 8'hed;
        my_rom[4837] = 8'hed;
        my_rom[4838] = 8'hed;
        my_rom[4839] = 8'he5;
        my_rom[4840] = 8'he5;
        my_rom[4841] = 8'he5;
        my_rom[4842] = 8'h93;
        my_rom[4843] = 8'h49;
        my_rom[4844] = 8'h53;
        my_rom[4845] = 8'h9b;
        my_rom[4846] = 8'h9b;
        my_rom[4847] = 8'h9b;
        my_rom[4848] = 8'h51;
        my_rom[4849] = 8'h49;
        my_rom[4850] = 8'h93;
        my_rom[4851] = 8'ha5;
        my_rom[4852] = 8'ha5;
        my_rom[4853] = 8'had;
        my_rom[4854] = 8'hef;
        my_rom[4855] = 8'hef;
        my_rom[4856] = 8'hef;
        my_rom[4857] = 8'hef;
        my_rom[4858] = 8'hef;
        my_rom[4859] = 8'hef;
        my_rom[4860] = 8'hef;
        my_rom[4861] = 8'hed;
        my_rom[4862] = 8'hed;
        my_rom[4863] = 8'hef;
        my_rom[4864] = 8'hef;
        my_rom[4865] = 8'haf;
        my_rom[4866] = 8'had;
        my_rom[4867] = 8'had;
        my_rom[4868] = 8'h8;
        my_rom[4869] = 8'h8;
        my_rom[4870] = 8'h8;
        my_rom[4871] = 8'ha;
        my_rom[4872] = 8'h8;
        my_rom[4873] = 8'h8;
        my_rom[4874] = 8'h8;
        my_rom[4875] = 8'h8;
        my_rom[4876] = 8'hf7;
        my_rom[4877] = 8'hf7;
        my_rom[4878] = 8'hf7;
        my_rom[4879] = 8'hf7;
        my_rom[4880] = 8'hf7;
        my_rom[4881] = 8'hf7;
        my_rom[4882] = 8'hf7;
        my_rom[4883] = 8'hf7;
        my_rom[4884] = 8'hf7;
        my_rom[4885] = 8'hf7;
        my_rom[4886] = 8'hf7;
        my_rom[4887] = 8'hf7;
        my_rom[4888] = 8'hf7;
        my_rom[4889] = 8'hf7;
        my_rom[4890] = 8'hf7;
        my_rom[4891] = 8'hf7;
        my_rom[4892] = 8'hf7;
        my_rom[4893] = 8'hf7;
        my_rom[4894] = 8'hef;
        my_rom[4895] = 8'hef;
        my_rom[4896] = 8'hed;
        my_rom[4897] = 8'hed;
        my_rom[4898] = 8'hed;
        my_rom[4899] = 8'hef;
        my_rom[4900] = 8'hef;
        my_rom[4901] = 8'he5;
        my_rom[4902] = 8'h9b;
        my_rom[4903] = 8'h9b;
        my_rom[4904] = 8'h9b;
        my_rom[4905] = 8'h9b;
        my_rom[4906] = 8'h9b;
        my_rom[4907] = 8'h9b;
        my_rom[4908] = 8'h9b;
        my_rom[4909] = 8'h9b;
        my_rom[4910] = 8'h9b;
        my_rom[4911] = 8'ha5;
        my_rom[4912] = 8'ha5;
        my_rom[4913] = 8'had;
        my_rom[4914] = 8'had;
        my_rom[4915] = 8'hef;
        my_rom[4916] = 8'hef;
        my_rom[4917] = 8'hef;
        my_rom[4918] = 8'hef;
        my_rom[4919] = 8'hed;
        my_rom[4920] = 8'hed;
        my_rom[4921] = 8'hed;
        my_rom[4922] = 8'hed;
        my_rom[4923] = 8'hef;
        my_rom[4924] = 8'hef;
        my_rom[4925] = 8'hef;
        my_rom[4926] = 8'had;
        my_rom[4927] = 8'hab;
        my_rom[4928] = 8'h8;
        my_rom[4929] = 8'h8;
        my_rom[4930] = 8'h8;
        my_rom[4931] = 8'ha;
        my_rom[4932] = 8'h8;
        my_rom[4933] = 8'h8;
        my_rom[4934] = 8'h8;
        my_rom[4935] = 8'h8;
        my_rom[4936] = 8'h8;
        my_rom[4937] = 8'hed;
        my_rom[4938] = 8'hed;
        my_rom[4939] = 8'hed;
        my_rom[4940] = 8'hed;
        my_rom[4941] = 8'hed;
        my_rom[4942] = 8'hed;
        my_rom[4943] = 8'hf7;
        my_rom[4944] = 8'hf7;
        my_rom[4945] = 8'hf7;
        my_rom[4946] = 8'hf7;
        my_rom[4947] = 8'hf7;
        my_rom[4948] = 8'hf7;
        my_rom[4949] = 8'hf7;
        my_rom[4950] = 8'hf7;
        my_rom[4951] = 8'hf7;
        my_rom[4952] = 8'hf7;
        my_rom[4953] = 8'hef;
        my_rom[4954] = 8'hed;
        my_rom[4955] = 8'hed;
        my_rom[4956] = 8'hed;
        my_rom[4957] = 8'hef;
        my_rom[4958] = 8'hef;
        my_rom[4959] = 8'hef;
        my_rom[4960] = 8'hef;
        my_rom[4961] = 8'hef;
        my_rom[4962] = 8'hed;
        my_rom[4963] = 8'he5;
        my_rom[4964] = 8'ha5;
        my_rom[4965] = 8'ha5;
        my_rom[4966] = 8'h9b;
        my_rom[4967] = 8'h9b;
        my_rom[4968] = 8'h9b;
        my_rom[4969] = 8'h9d;
        my_rom[4970] = 8'ha5;
        my_rom[4971] = 8'ha5;
        my_rom[4972] = 8'had;
        my_rom[4973] = 8'had;
        my_rom[4974] = 8'hed;
        my_rom[4975] = 8'hed;
        my_rom[4976] = 8'hed;
        my_rom[4977] = 8'hed;
        my_rom[4978] = 8'hed;
        my_rom[4979] = 8'hed;
        my_rom[4980] = 8'hed;
        my_rom[4981] = 8'hed;
        my_rom[4982] = 8'hed;
        my_rom[4983] = 8'hed;
        my_rom[4984] = 8'hed;
        my_rom[4985] = 8'hed;
        my_rom[4986] = 8'had;
        my_rom[4987] = 8'h8;
        my_rom[4988] = 8'h8;
        my_rom[4989] = 8'h8;
        my_rom[4990] = 8'h8;
        my_rom[4991] = 8'ha;
        my_rom[4992] = 8'h8;
        my_rom[4993] = 8'h8;
        my_rom[4994] = 8'h8;
        my_rom[4995] = 8'h8;
        my_rom[4996] = 8'h8;
        my_rom[4997] = 8'h8;
        my_rom[4998] = 8'h8;
        my_rom[4999] = 8'h8;
        my_rom[5000] = 8'ha5;
        my_rom[5001] = 8'ha3;
        my_rom[5002] = 8'ha5;
        my_rom[5003] = 8'hf7;
        my_rom[5004] = 8'hf7;
        my_rom[5005] = 8'hf7;
        my_rom[5006] = 8'hf7;
        my_rom[5007] = 8'hf7;
        my_rom[5008] = 8'hf7;
        my_rom[5009] = 8'hf7;
        my_rom[5010] = 8'hf7;
        my_rom[5011] = 8'hf7;
        my_rom[5012] = 8'hf7;
        my_rom[5013] = 8'hed;
        my_rom[5014] = 8'hed;
        my_rom[5015] = 8'hed;
        my_rom[5016] = 8'hef;
        my_rom[5017] = 8'hf7;
        my_rom[5018] = 8'hf7;
        my_rom[5019] = 8'hf7;
        my_rom[5020] = 8'hf7;
        my_rom[5021] = 8'hef;
        my_rom[5022] = 8'hef;
        my_rom[5023] = 8'hef;
        my_rom[5024] = 8'hed;
        my_rom[5025] = 8'ha5;
        my_rom[5026] = 8'ha5;
        my_rom[5027] = 8'ha5;
        my_rom[5028] = 8'ha5;
        my_rom[5029] = 8'ha5;
        my_rom[5030] = 8'ha5;
        my_rom[5031] = 8'ha5;
        my_rom[5032] = 8'haf;
        my_rom[5033] = 8'hef;
        my_rom[5034] = 8'hed;
        my_rom[5035] = 8'hed;
        my_rom[5036] = 8'hed;
        my_rom[5037] = 8'hed;
        my_rom[5038] = 8'hed;
        my_rom[5039] = 8'hed;
        my_rom[5040] = 8'hed;
        my_rom[5041] = 8'hed;
        my_rom[5042] = 8'had;
        my_rom[5043] = 8'ha5;
        my_rom[5044] = 8'ha5;
        my_rom[5045] = 8'h8;
        my_rom[5046] = 8'h8;
        my_rom[5047] = 8'h8;
        my_rom[5048] = 8'h8;
        my_rom[5049] = 8'h8;
        my_rom[5050] = 8'h8;
        my_rom[5051] = 8'ha;
        my_rom[5052] = 8'h8;
        my_rom[5053] = 8'h8;
        my_rom[5054] = 8'h8;
        my_rom[5055] = 8'h8;
        my_rom[5056] = 8'h8;
        my_rom[5057] = 8'h8;
        my_rom[5058] = 8'h8;
        my_rom[5059] = 8'h8;
        my_rom[5060] = 8'h8;
        my_rom[5061] = 8'h8;
        my_rom[5062] = 8'ha5;
        my_rom[5063] = 8'hf7;
        my_rom[5064] = 8'hf7;
        my_rom[5065] = 8'hf7;
        my_rom[5066] = 8'hf7;
        my_rom[5067] = 8'hf7;
        my_rom[5068] = 8'hf7;
        my_rom[5069] = 8'hf7;
        my_rom[5070] = 8'hf7;
        my_rom[5071] = 8'hf7;
        my_rom[5072] = 8'hed;
        my_rom[5073] = 8'hed;
        my_rom[5074] = 8'hed;
        my_rom[5075] = 8'hef;
        my_rom[5076] = 8'hf7;
        my_rom[5077] = 8'hf7;
        my_rom[5078] = 8'hf7;
        my_rom[5079] = 8'hf7;
        my_rom[5080] = 8'hf7;
        my_rom[5081] = 8'hef;
        my_rom[5082] = 8'hef;
        my_rom[5083] = 8'hef;
        my_rom[5084] = 8'hed;
        my_rom[5085] = 8'ha5;
        my_rom[5086] = 8'ha5;
        my_rom[5087] = 8'ha5;
        my_rom[5088] = 8'ha5;
        my_rom[5089] = 8'ha5;
        my_rom[5090] = 8'ha5;
        my_rom[5091] = 8'haf;
        my_rom[5092] = 8'haf;
        my_rom[5093] = 8'hef;
        my_rom[5094] = 8'hed;
        my_rom[5095] = 8'hed;
        my_rom[5096] = 8'hed;
        my_rom[5097] = 8'hed;
        my_rom[5098] = 8'hed;
        my_rom[5099] = 8'hed;
        my_rom[5100] = 8'hed;
        my_rom[5101] = 8'hed;
        my_rom[5102] = 8'ha5;
        my_rom[5103] = 8'h8;
        my_rom[5104] = 8'h8;
        my_rom[5105] = 8'h8;
        my_rom[5106] = 8'h8;
        my_rom[5107] = 8'h8;
        my_rom[5108] = 8'h8;
        my_rom[5109] = 8'h8;
        my_rom[5110] = 8'h8;
        my_rom[5111] = 8'ha;
        my_rom[5112] = 8'h8;
        my_rom[5113] = 8'h8;
        my_rom[5114] = 8'h8;
        my_rom[5115] = 8'h8;
        my_rom[5116] = 8'h8;
        my_rom[5117] = 8'h8;
        my_rom[5118] = 8'h8;
        my_rom[5119] = 8'h8;
        my_rom[5120] = 8'h8;
        my_rom[5121] = 8'h8;
        my_rom[5122] = 8'ha5;
        my_rom[5123] = 8'hf7;
        my_rom[5124] = 8'hf7;
        my_rom[5125] = 8'hf7;
        my_rom[5126] = 8'hf7;
        my_rom[5127] = 8'hf7;
        my_rom[5128] = 8'hf7;
        my_rom[5129] = 8'hf7;
        my_rom[5130] = 8'hf7;
        my_rom[5131] = 8'hf7;
        my_rom[5132] = 8'hed;
        my_rom[5133] = 8'hed;
        my_rom[5134] = 8'hef;
        my_rom[5135] = 8'hef;
        my_rom[5136] = 8'hef;
        my_rom[5137] = 8'hf7;
        my_rom[5138] = 8'hf7;
        my_rom[5139] = 8'hf7;
        my_rom[5140] = 8'hf7;
        my_rom[5141] = 8'hf7;
        my_rom[5142] = 8'hef;
        my_rom[5143] = 8'hef;
        my_rom[5144] = 8'hef;
        my_rom[5145] = 8'hef;
        my_rom[5146] = 8'he5;
        my_rom[5147] = 8'hed;
        my_rom[5148] = 8'ha5;
        my_rom[5149] = 8'ha5;
        my_rom[5150] = 8'had;
        my_rom[5151] = 8'had;
        my_rom[5152] = 8'had;
        my_rom[5153] = 8'had;
        my_rom[5154] = 8'hed;
        my_rom[5155] = 8'hed;
        my_rom[5156] = 8'hed;
        my_rom[5157] = 8'hed;
        my_rom[5158] = 8'hed;
        my_rom[5159] = 8'hed;
        my_rom[5160] = 8'hed;
        my_rom[5161] = 8'hed;
        my_rom[5162] = 8'ha5;
        my_rom[5163] = 8'h8;
        my_rom[5164] = 8'h8;
        my_rom[5165] = 8'h8;
        my_rom[5166] = 8'h8;
        my_rom[5167] = 8'h8;
        my_rom[5168] = 8'h8;
        my_rom[5169] = 8'h8;
        my_rom[5170] = 8'h8;
        my_rom[5171] = 8'ha;
        my_rom[5172] = 8'h8;
        my_rom[5173] = 8'h8;
        my_rom[5174] = 8'h8;
        my_rom[5175] = 8'h8;
        my_rom[5176] = 8'h8;
        my_rom[5177] = 8'h8;
        my_rom[5178] = 8'h8;
        my_rom[5179] = 8'h8;
        my_rom[5180] = 8'h8;
        my_rom[5181] = 8'h8;
        my_rom[5182] = 8'had;
        my_rom[5183] = 8'hf7;
        my_rom[5184] = 8'hf7;
        my_rom[5185] = 8'hf7;
        my_rom[5186] = 8'hf7;
        my_rom[5187] = 8'hf7;
        my_rom[5188] = 8'hf7;
        my_rom[5189] = 8'hf7;
        my_rom[5190] = 8'hf7;
        my_rom[5191] = 8'hed;
        my_rom[5192] = 8'hed;
        my_rom[5193] = 8'hed;
        my_rom[5194] = 8'hed;
        my_rom[5195] = 8'hed;
        my_rom[5196] = 8'hed;
        my_rom[5197] = 8'hef;
        my_rom[5198] = 8'hef;
        my_rom[5199] = 8'hef;
        my_rom[5200] = 8'hef;
        my_rom[5201] = 8'hef;
        my_rom[5202] = 8'hef;
        my_rom[5203] = 8'hef;
        my_rom[5204] = 8'hef;
        my_rom[5205] = 8'hef;
        my_rom[5206] = 8'hef;
        my_rom[5207] = 8'he5;
        my_rom[5208] = 8'had;
        my_rom[5209] = 8'had;
        my_rom[5210] = 8'had;
        my_rom[5211] = 8'had;
        my_rom[5212] = 8'had;
        my_rom[5213] = 8'ha5;
        my_rom[5214] = 8'ha5;
        my_rom[5215] = 8'he5;
        my_rom[5216] = 8'hed;
        my_rom[5217] = 8'hed;
        my_rom[5218] = 8'he5;
        my_rom[5219] = 8'ha5;
        my_rom[5220] = 8'had;
        my_rom[5221] = 8'hed;
        my_rom[5222] = 8'ha5;
        my_rom[5223] = 8'h8;
        my_rom[5224] = 8'h8;
        my_rom[5225] = 8'h8;
        my_rom[5226] = 8'h8;
        my_rom[5227] = 8'h8;
        my_rom[5228] = 8'h8;
        my_rom[5229] = 8'h8;
        my_rom[5230] = 8'h8;
        my_rom[5231] = 8'ha;
        my_rom[5232] = 8'h8;
        my_rom[5233] = 8'h8;
        my_rom[5234] = 8'h8;
        my_rom[5235] = 8'h8;
        my_rom[5236] = 8'h8;
        my_rom[5237] = 8'h8;
        my_rom[5238] = 8'h8;
        my_rom[5239] = 8'h8;
        my_rom[5240] = 8'h8;
        my_rom[5241] = 8'h8;
        my_rom[5242] = 8'ha5;
        my_rom[5243] = 8'hf5;
        my_rom[5244] = 8'hf7;
        my_rom[5245] = 8'hf7;
        my_rom[5246] = 8'hf7;
        my_rom[5247] = 8'hf7;
        my_rom[5248] = 8'hf7;
        my_rom[5249] = 8'hf7;
        my_rom[5250] = 8'hf5;
        my_rom[5251] = 8'hed;
        my_rom[5252] = 8'hed;
        my_rom[5253] = 8'hed;
        my_rom[5254] = 8'hed;
        my_rom[5255] = 8'hed;
        my_rom[5256] = 8'hed;
        my_rom[5257] = 8'hed;
        my_rom[5258] = 8'hef;
        my_rom[5259] = 8'hef;
        my_rom[5260] = 8'hef;
        my_rom[5261] = 8'hed;
        my_rom[5262] = 8'he5;
        my_rom[5263] = 8'ha5;
        my_rom[5264] = 8'h9b;
        my_rom[5265] = 8'h9d;
        my_rom[5266] = 8'h9b;
        my_rom[5267] = 8'h9b;
        my_rom[5268] = 8'h9d;
        my_rom[5269] = 8'ha5;
        my_rom[5270] = 8'ha5;
        my_rom[5271] = 8'had;
        my_rom[5272] = 8'ha5;
        my_rom[5273] = 8'ha5;
        my_rom[5274] = 8'ha5;
        my_rom[5275] = 8'ha5;
        my_rom[5276] = 8'ha5;
        my_rom[5277] = 8'had;
        my_rom[5278] = 8'ha5;
        my_rom[5279] = 8'had;
        my_rom[5280] = 8'had;
        my_rom[5281] = 8'hed;
        my_rom[5282] = 8'ha5;
        my_rom[5283] = 8'h8;
        my_rom[5284] = 8'h8;
        my_rom[5285] = 8'h8;
        my_rom[5286] = 8'h8;
        my_rom[5287] = 8'h8;
        my_rom[5288] = 8'h8;
        my_rom[5289] = 8'h8;
        my_rom[5290] = 8'h8;
        my_rom[5291] = 8'ha;
        my_rom[5292] = 8'h8;
        my_rom[5293] = 8'h8;
        my_rom[5294] = 8'h8;
        my_rom[5295] = 8'h8;
        my_rom[5296] = 8'h8;
        my_rom[5297] = 8'h8;
        my_rom[5298] = 8'h8;
        my_rom[5299] = 8'h8;
        my_rom[5300] = 8'h8;
        my_rom[5301] = 8'h8;
        my_rom[5302] = 8'ha5;
        my_rom[5303] = 8'hed;
        my_rom[5304] = 8'hf7;
        my_rom[5305] = 8'hf7;
        my_rom[5306] = 8'hf7;
        my_rom[5307] = 8'hf7;
        my_rom[5308] = 8'hf7;
        my_rom[5309] = 8'hf7;
        my_rom[5310] = 8'hf5;
        my_rom[5311] = 8'hed;
        my_rom[5312] = 8'hed;
        my_rom[5313] = 8'hed;
        my_rom[5314] = 8'hed;
        my_rom[5315] = 8'ha5;
        my_rom[5316] = 8'ha5;
        my_rom[5317] = 8'ha5;
        my_rom[5318] = 8'ha5;
        my_rom[5319] = 8'ha5;
        my_rom[5320] = 8'h9b;
        my_rom[5321] = 8'h9b;
        my_rom[5322] = 8'h93;
        my_rom[5323] = 8'h93;
        my_rom[5324] = 8'h93;
        my_rom[5325] = 8'h93;
        my_rom[5326] = 8'h93;
        my_rom[5327] = 8'h93;
        my_rom[5328] = 8'h93;
        my_rom[5329] = 8'h93;
        my_rom[5330] = 8'h9b;
        my_rom[5331] = 8'h9d;
        my_rom[5332] = 8'ha5;
        my_rom[5333] = 8'ha5;
        my_rom[5334] = 8'ha5;
        my_rom[5335] = 8'ha5;
        my_rom[5336] = 8'ha5;
        my_rom[5337] = 8'ha5;
        my_rom[5338] = 8'ha5;
        my_rom[5339] = 8'had;
        my_rom[5340] = 8'had;
        my_rom[5341] = 8'had;
        my_rom[5342] = 8'h5b;
        my_rom[5343] = 8'h8;
        my_rom[5344] = 8'h8;
        my_rom[5345] = 8'h8;
        my_rom[5346] = 8'h8;
        my_rom[5347] = 8'h8;
        my_rom[5348] = 8'h8;
        my_rom[5349] = 8'h8;
        my_rom[5350] = 8'h8;
        my_rom[5351] = 8'ha;
        my_rom[5352] = 8'h8;
        my_rom[5353] = 8'h8;
        my_rom[5354] = 8'h8;
        my_rom[5355] = 8'h8;
        my_rom[5356] = 8'h8;
        my_rom[5357] = 8'h8;
        my_rom[5358] = 8'h8;
        my_rom[5359] = 8'h8;
        my_rom[5360] = 8'h8;
        my_rom[5361] = 8'h8;
        my_rom[5362] = 8'ha5;
        my_rom[5363] = 8'hed;
        my_rom[5364] = 8'hf7;
        my_rom[5365] = 8'hf7;
        my_rom[5366] = 8'hf7;
        my_rom[5367] = 8'hf7;
        my_rom[5368] = 8'hf7;
        my_rom[5369] = 8'hed;
        my_rom[5370] = 8'hed;
        my_rom[5371] = 8'hed;
        my_rom[5372] = 8'hed;
        my_rom[5373] = 8'hed;
        my_rom[5374] = 8'ha5;
        my_rom[5375] = 8'ha5;
        my_rom[5376] = 8'h9b;
        my_rom[5377] = 8'h93;
        my_rom[5378] = 8'h53;
        my_rom[5379] = 8'h53;
        my_rom[5380] = 8'h93;
        my_rom[5381] = 8'h93;
        my_rom[5382] = 8'h93;
        my_rom[5383] = 8'h93;
        my_rom[5384] = 8'h93;
        my_rom[5385] = 8'h8b;
        my_rom[5386] = 8'h4b;
        my_rom[5387] = 8'h4b;
        my_rom[5388] = 8'h4b;
        my_rom[5389] = 8'h53;
        my_rom[5390] = 8'h53;
        my_rom[5391] = 8'h53;
        my_rom[5392] = 8'h53;
        my_rom[5393] = 8'h9b;
        my_rom[5394] = 8'h9b;
        my_rom[5395] = 8'ha5;
        my_rom[5396] = 8'ha5;
        my_rom[5397] = 8'ha5;
        my_rom[5398] = 8'ha5;
        my_rom[5399] = 8'ha5;
        my_rom[5400] = 8'had;
        my_rom[5401] = 8'had;
        my_rom[5402] = 8'h8;
        my_rom[5403] = 8'h8;
        my_rom[5404] = 8'h8;
        my_rom[5405] = 8'h8;
        my_rom[5406] = 8'h8;
        my_rom[5407] = 8'h8;
        my_rom[5408] = 8'h8;
        my_rom[5409] = 8'h8;
        my_rom[5410] = 8'h8;
        my_rom[5411] = 8'ha;
        my_rom[5412] = 8'h8;
        my_rom[5413] = 8'h8;
        my_rom[5414] = 8'h8;
        my_rom[5415] = 8'h8;
        my_rom[5416] = 8'h8;
        my_rom[5417] = 8'h8;
        my_rom[5418] = 8'h8;
        my_rom[5419] = 8'h8;
        my_rom[5420] = 8'h8;
        my_rom[5421] = 8'h8;
        my_rom[5422] = 8'h8;
        my_rom[5423] = 8'had;
        my_rom[5424] = 8'hf7;
        my_rom[5425] = 8'hf5;
        my_rom[5426] = 8'hf7;
        my_rom[5427] = 8'hf7;
        my_rom[5428] = 8'hf7;
        my_rom[5429] = 8'hed;
        my_rom[5430] = 8'hed;
        my_rom[5431] = 8'hed;
        my_rom[5432] = 8'hed;
        my_rom[5433] = 8'hed;
        my_rom[5434] = 8'ha5;
        my_rom[5435] = 8'h9b;
        my_rom[5436] = 8'h9b;
        my_rom[5437] = 8'ha5;
        my_rom[5438] = 8'h9d;
        my_rom[5439] = 8'h9d;
        my_rom[5440] = 8'he5;
        my_rom[5441] = 8'he7;
        my_rom[5442] = 8'hef;
        my_rom[5443] = 8'hef;
        my_rom[5444] = 8'he7;
        my_rom[5445] = 8'he5;
        my_rom[5446] = 8'ha5;
        my_rom[5447] = 8'h9d;
        my_rom[5448] = 8'h9d;
        my_rom[5449] = 8'h9d;
        my_rom[5450] = 8'h9d;
        my_rom[5451] = 8'h53;
        my_rom[5452] = 8'h53;
        my_rom[5453] = 8'h93;
        my_rom[5454] = 8'h9b;
        my_rom[5455] = 8'ha5;
        my_rom[5456] = 8'ha5;
        my_rom[5457] = 8'ha5;
        my_rom[5458] = 8'ha5;
        my_rom[5459] = 8'had;
        my_rom[5460] = 8'hed;
        my_rom[5461] = 8'had;
        my_rom[5462] = 8'h8;
        my_rom[5463] = 8'h8;
        my_rom[5464] = 8'h8;
        my_rom[5465] = 8'h8;
        my_rom[5466] = 8'h8;
        my_rom[5467] = 8'h8;
        my_rom[5468] = 8'h8;
        my_rom[5469] = 8'h8;
        my_rom[5470] = 8'h8;
        my_rom[5471] = 8'ha;
        my_rom[5472] = 8'h8;
        my_rom[5473] = 8'h8;
        my_rom[5474] = 8'h8;
        my_rom[5475] = 8'h8;
        my_rom[5476] = 8'h8;
        my_rom[5477] = 8'h8;
        my_rom[5478] = 8'h8;
        my_rom[5479] = 8'h8;
        my_rom[5480] = 8'h8;
        my_rom[5481] = 8'h8;
        my_rom[5482] = 8'h8;
        my_rom[5483] = 8'had;
        my_rom[5484] = 8'hf7;
        my_rom[5485] = 8'hf5;
        my_rom[5486] = 8'hf5;
        my_rom[5487] = 8'hf5;
        my_rom[5488] = 8'hed;
        my_rom[5489] = 8'hed;
        my_rom[5490] = 8'hed;
        my_rom[5491] = 8'hed;
        my_rom[5492] = 8'hed;
        my_rom[5493] = 8'hed;
        my_rom[5494] = 8'ha5;
        my_rom[5495] = 8'ha5;
        my_rom[5496] = 8'ha5;
        my_rom[5497] = 8'hed;
        my_rom[5498] = 8'hed;
        my_rom[5499] = 8'hed;
        my_rom[5500] = 8'he5;
        my_rom[5501] = 8'he5;
        my_rom[5502] = 8'he5;
        my_rom[5503] = 8'he7;
        my_rom[5504] = 8'he5;
        my_rom[5505] = 8'he5;
        my_rom[5506] = 8'he5;
        my_rom[5507] = 8'ha5;
        my_rom[5508] = 8'h9d;
        my_rom[5509] = 8'h9d;
        my_rom[5510] = 8'h9d;
        my_rom[5511] = 8'h9d;
        my_rom[5512] = 8'ha5;
        my_rom[5513] = 8'ha5;
        my_rom[5514] = 8'h9b;
        my_rom[5515] = 8'ha5;
        my_rom[5516] = 8'ha5;
        my_rom[5517] = 8'ha5;
        my_rom[5518] = 8'ha5;
        my_rom[5519] = 8'had;
        my_rom[5520] = 8'had;
        my_rom[5521] = 8'ha5;
        my_rom[5522] = 8'h8;
        my_rom[5523] = 8'h8;
        my_rom[5524] = 8'h8;
        my_rom[5525] = 8'h8;
        my_rom[5526] = 8'h8;
        my_rom[5527] = 8'h8;
        my_rom[5528] = 8'h8;
        my_rom[5529] = 8'h8;
        my_rom[5530] = 8'h8;
        my_rom[5531] = 8'ha;
        my_rom[5532] = 8'h8;
        my_rom[5533] = 8'h8;
        my_rom[5534] = 8'h8;
        my_rom[5535] = 8'h8;
        my_rom[5536] = 8'h8;
        my_rom[5537] = 8'h8;
        my_rom[5538] = 8'h8;
        my_rom[5539] = 8'h8;
        my_rom[5540] = 8'h8;
        my_rom[5541] = 8'h8;
        my_rom[5542] = 8'h8;
        my_rom[5543] = 8'had;
        my_rom[5544] = 8'hf7;
        my_rom[5545] = 8'hf5;
        my_rom[5546] = 8'hf5;
        my_rom[5547] = 8'hed;
        my_rom[5548] = 8'hed;
        my_rom[5549] = 8'hed;
        my_rom[5550] = 8'hed;
        my_rom[5551] = 8'hed;
        my_rom[5552] = 8'hed;
        my_rom[5553] = 8'hed;
        my_rom[5554] = 8'ha5;
        my_rom[5555] = 8'ha5;
        my_rom[5556] = 8'hed;
        my_rom[5557] = 8'hed;
        my_rom[5558] = 8'hed;
        my_rom[5559] = 8'hed;
        my_rom[5560] = 8'hed;
        my_rom[5561] = 8'he5;
        my_rom[5562] = 8'hdd;
        my_rom[5563] = 8'h9d;
        my_rom[5564] = 8'h9d;
        my_rom[5565] = 8'h9d;
        my_rom[5566] = 8'h9d;
        my_rom[5567] = 8'h9d;
        my_rom[5568] = 8'h9d;
        my_rom[5569] = 8'h9d;
        my_rom[5570] = 8'h9d;
        my_rom[5571] = 8'ha5;
        my_rom[5572] = 8'ha5;
        my_rom[5573] = 8'ha5;
        my_rom[5574] = 8'ha5;
        my_rom[5575] = 8'ha5;
        my_rom[5576] = 8'ha5;
        my_rom[5577] = 8'ha5;
        my_rom[5578] = 8'ha5;
        my_rom[5579] = 8'had;
        my_rom[5580] = 8'ha5;
        my_rom[5581] = 8'h53;
        my_rom[5582] = 8'h8;
        my_rom[5583] = 8'h8;
        my_rom[5584] = 8'h8;
        my_rom[5585] = 8'h8;
        my_rom[5586] = 8'h8;
        my_rom[5587] = 8'h8;
        my_rom[5588] = 8'h8;
        my_rom[5589] = 8'h8;
        my_rom[5590] = 8'h8;
        my_rom[5591] = 8'ha;
        my_rom[5592] = 8'h8;
        my_rom[5593] = 8'h8;
        my_rom[5594] = 8'h8;
        my_rom[5595] = 8'h8;
        my_rom[5596] = 8'h8;
        my_rom[5597] = 8'h8;
        my_rom[5598] = 8'h8;
        my_rom[5599] = 8'h8;
        my_rom[5600] = 8'h8;
        my_rom[5601] = 8'h8;
        my_rom[5602] = 8'h8;
        my_rom[5603] = 8'had;
        my_rom[5604] = 8'hf7;
        my_rom[5605] = 8'hf5;
        my_rom[5606] = 8'hed;
        my_rom[5607] = 8'hed;
        my_rom[5608] = 8'hed;
        my_rom[5609] = 8'hed;
        my_rom[5610] = 8'hed;
        my_rom[5611] = 8'hed;
        my_rom[5612] = 8'hed;
        my_rom[5613] = 8'hed;
        my_rom[5614] = 8'hed;
        my_rom[5615] = 8'hed;
        my_rom[5616] = 8'hed;
        my_rom[5617] = 8'hed;
        my_rom[5618] = 8'hed;
        my_rom[5619] = 8'hed;
        my_rom[5620] = 8'hed;
        my_rom[5621] = 8'ha5;
        my_rom[5622] = 8'h9b;
        my_rom[5623] = 8'h9b;
        my_rom[5624] = 8'h9b;
        my_rom[5625] = 8'h9b;
        my_rom[5626] = 8'h93;
        my_rom[5627] = 8'h93;
        my_rom[5628] = 8'h9b;
        my_rom[5629] = 8'h9b;
        my_rom[5630] = 8'ha5;
        my_rom[5631] = 8'ha5;
        my_rom[5632] = 8'ha5;
        my_rom[5633] = 8'ha5;
        my_rom[5634] = 8'ha5;
        my_rom[5635] = 8'ha5;
        my_rom[5636] = 8'ha5;
        my_rom[5637] = 8'ha5;
        my_rom[5638] = 8'ha5;
        my_rom[5639] = 8'had;
        my_rom[5640] = 8'h5b;
        my_rom[5641] = 8'h8;
        my_rom[5642] = 8'h8;
        my_rom[5643] = 8'h8;
        my_rom[5644] = 8'h8;
        my_rom[5645] = 8'h8;
        my_rom[5646] = 8'h8;
        my_rom[5647] = 8'h8;
        my_rom[5648] = 8'h8;
        my_rom[5649] = 8'h8;
        my_rom[5650] = 8'h8;
        my_rom[5651] = 8'ha;
        my_rom[5652] = 8'h8;
        my_rom[5653] = 8'h8;
        my_rom[5654] = 8'h8;
        my_rom[5655] = 8'h8;
        my_rom[5656] = 8'h8;
        my_rom[5657] = 8'h8;
        my_rom[5658] = 8'h8;
        my_rom[5659] = 8'h8;
        my_rom[5660] = 8'h8;
        my_rom[5661] = 8'h8;
        my_rom[5662] = 8'h8;
        my_rom[5663] = 8'had;
        my_rom[5664] = 8'hf7;
        my_rom[5665] = 8'hf7;
        my_rom[5666] = 8'hed;
        my_rom[5667] = 8'hed;
        my_rom[5668] = 8'hed;
        my_rom[5669] = 8'hed;
        my_rom[5670] = 8'hed;
        my_rom[5671] = 8'hed;
        my_rom[5672] = 8'hed;
        my_rom[5673] = 8'hed;
        my_rom[5674] = 8'hed;
        my_rom[5675] = 8'hed;
        my_rom[5676] = 8'hed;
        my_rom[5677] = 8'hed;
        my_rom[5678] = 8'hed;
        my_rom[5679] = 8'hed;
        my_rom[5680] = 8'he5;
        my_rom[5681] = 8'ha5;
        my_rom[5682] = 8'ha3;
        my_rom[5683] = 8'h9b;
        my_rom[5684] = 8'h9b;
        my_rom[5685] = 8'h9b;
        my_rom[5686] = 8'h9b;
        my_rom[5687] = 8'h9b;
        my_rom[5688] = 8'h9b;
        my_rom[5689] = 8'h9b;
        my_rom[5690] = 8'ha3;
        my_rom[5691] = 8'ha5;
        my_rom[5692] = 8'ha5;
        my_rom[5693] = 8'ha5;
        my_rom[5694] = 8'ha5;
        my_rom[5695] = 8'ha5;
        my_rom[5696] = 8'ha5;
        my_rom[5697] = 8'ha5;
        my_rom[5698] = 8'had;
        my_rom[5699] = 8'ha5;
        my_rom[5700] = 8'h53;
        my_rom[5701] = 8'h8;
        my_rom[5702] = 8'h8;
        my_rom[5703] = 8'h8;
        my_rom[5704] = 8'h8;
        my_rom[5705] = 8'h8;
        my_rom[5706] = 8'h8;
        my_rom[5707] = 8'h8;
        my_rom[5708] = 8'h8;
        my_rom[5709] = 8'h8;
        my_rom[5710] = 8'h8;
        my_rom[5711] = 8'ha;
        my_rom[5712] = 8'h8;
        my_rom[5713] = 8'h8;
        my_rom[5714] = 8'h8;
        my_rom[5715] = 8'h8;
        my_rom[5716] = 8'h8;
        my_rom[5717] = 8'h8;
        my_rom[5718] = 8'h8;
        my_rom[5719] = 8'h8;
        my_rom[5720] = 8'h8;
        my_rom[5721] = 8'h8;
        my_rom[5722] = 8'h8;
        my_rom[5723] = 8'had;
        my_rom[5724] = 8'hf7;
        my_rom[5725] = 8'hf7;
        my_rom[5726] = 8'hed;
        my_rom[5727] = 8'hed;
        my_rom[5728] = 8'hed;
        my_rom[5729] = 8'hed;
        my_rom[5730] = 8'hed;
        my_rom[5731] = 8'hed;
        my_rom[5732] = 8'hed;
        my_rom[5733] = 8'hed;
        my_rom[5734] = 8'hed;
        my_rom[5735] = 8'hed;
        my_rom[5736] = 8'hed;
        my_rom[5737] = 8'hed;
        my_rom[5738] = 8'hed;
        my_rom[5739] = 8'hed;
        my_rom[5740] = 8'he5;
        my_rom[5741] = 8'ha5;
        my_rom[5742] = 8'ha3;
        my_rom[5743] = 8'h9b;
        my_rom[5744] = 8'h9b;
        my_rom[5745] = 8'h9b;
        my_rom[5746] = 8'h9b;
        my_rom[5747] = 8'h9b;
        my_rom[5748] = 8'h9b;
        my_rom[5749] = 8'h9b;
        my_rom[5750] = 8'ha3;
        my_rom[5751] = 8'ha5;
        my_rom[5752] = 8'ha5;
        my_rom[5753] = 8'ha5;
        my_rom[5754] = 8'ha5;
        my_rom[5755] = 8'ha5;
        my_rom[5756] = 8'ha5;
        my_rom[5757] = 8'ha5;
        my_rom[5758] = 8'ha5;
        my_rom[5759] = 8'h5b;
        my_rom[5760] = 8'h53;
        my_rom[5761] = 8'h8;
        my_rom[5762] = 8'h8;
        my_rom[5763] = 8'h8;
        my_rom[5764] = 8'h8;
        my_rom[5765] = 8'h8;
        my_rom[5766] = 8'h8;
        my_rom[5767] = 8'h8;
        my_rom[5768] = 8'h8;
        my_rom[5769] = 8'h8;
        my_rom[5770] = 8'h8;
        my_rom[5771] = 8'ha;
        my_rom[5772] = 8'h8;
        my_rom[5773] = 8'h8;
        my_rom[5774] = 8'h8;
        my_rom[5775] = 8'h8;
        my_rom[5776] = 8'h8;
        my_rom[5777] = 8'h8;
        my_rom[5778] = 8'h8;
        my_rom[5779] = 8'h8;
        my_rom[5780] = 8'h8;
        my_rom[5781] = 8'h8;
        my_rom[5782] = 8'h8;
        my_rom[5783] = 8'hff;
        my_rom[5784] = 8'hf7;
        my_rom[5785] = 8'hf7;
        my_rom[5786] = 8'hf7;
        my_rom[5787] = 8'hed;
        my_rom[5788] = 8'hed;
        my_rom[5789] = 8'hed;
        my_rom[5790] = 8'hed;
        my_rom[5791] = 8'hed;
        my_rom[5792] = 8'hed;
        my_rom[5793] = 8'hed;
        my_rom[5794] = 8'hed;
        my_rom[5795] = 8'hed;
        my_rom[5796] = 8'hed;
        my_rom[5797] = 8'hed;
        my_rom[5798] = 8'hed;
        my_rom[5799] = 8'hed;
        my_rom[5800] = 8'he5;
        my_rom[5801] = 8'ha5;
        my_rom[5802] = 8'h9b;
        my_rom[5803] = 8'h9b;
        my_rom[5804] = 8'h9b;
        my_rom[5805] = 8'h9b;
        my_rom[5806] = 8'h9b;
        my_rom[5807] = 8'h9b;
        my_rom[5808] = 8'h9b;
        my_rom[5809] = 8'h9b;
        my_rom[5810] = 8'ha5;
        my_rom[5811] = 8'ha5;
        my_rom[5812] = 8'ha5;
        my_rom[5813] = 8'ha5;
        my_rom[5814] = 8'ha5;
        my_rom[5815] = 8'ha5;
        my_rom[5816] = 8'ha5;
        my_rom[5817] = 8'ha5;
        my_rom[5818] = 8'h9b;
        my_rom[5819] = 8'h53;
        my_rom[5820] = 8'h8;
        my_rom[5821] = 8'h8;
        my_rom[5822] = 8'h8;
        my_rom[5823] = 8'h8;
        my_rom[5824] = 8'h8;
        my_rom[5825] = 8'h8;
        my_rom[5826] = 8'h8;
        my_rom[5827] = 8'h8;
        my_rom[5828] = 8'h8;
        my_rom[5829] = 8'h8;
        my_rom[5830] = 8'h8;
        my_rom[5831] = 8'ha;
        my_rom[5832] = 8'h8;
        my_rom[5833] = 8'h8;
        my_rom[5834] = 8'h8;
        my_rom[5835] = 8'h8;
        my_rom[5836] = 8'h8;
        my_rom[5837] = 8'h8;
        my_rom[5838] = 8'h8;
        my_rom[5839] = 8'h8;
        my_rom[5840] = 8'h8;
        my_rom[5841] = 8'h8;
        my_rom[5842] = 8'h8;
        my_rom[5843] = 8'hf7;
        my_rom[5844] = 8'hf7;
        my_rom[5845] = 8'hf7;
        my_rom[5846] = 8'hf7;
        my_rom[5847] = 8'hf5;
        my_rom[5848] = 8'hed;
        my_rom[5849] = 8'hed;
        my_rom[5850] = 8'hed;
        my_rom[5851] = 8'hed;
        my_rom[5852] = 8'hed;
        my_rom[5853] = 8'hed;
        my_rom[5854] = 8'hed;
        my_rom[5855] = 8'hed;
        my_rom[5856] = 8'hed;
        my_rom[5857] = 8'hed;
        my_rom[5858] = 8'hed;
        my_rom[5859] = 8'hed;
        my_rom[5860] = 8'hed;
        my_rom[5861] = 8'he5;
        my_rom[5862] = 8'ha5;
        my_rom[5863] = 8'ha5;
        my_rom[5864] = 8'ha5;
        my_rom[5865] = 8'ha5;
        my_rom[5866] = 8'ha5;
        my_rom[5867] = 8'ha5;
        my_rom[5868] = 8'ha5;
        my_rom[5869] = 8'ha5;
        my_rom[5870] = 8'ha5;
        my_rom[5871] = 8'ha5;
        my_rom[5872] = 8'ha5;
        my_rom[5873] = 8'ha5;
        my_rom[5874] = 8'ha5;
        my_rom[5875] = 8'ha5;
        my_rom[5876] = 8'ha5;
        my_rom[5877] = 8'ha5;
        my_rom[5878] = 8'h53;
        my_rom[5879] = 8'h8;
        my_rom[5880] = 8'h8;
        my_rom[5881] = 8'h8;
        my_rom[5882] = 8'h8;
        my_rom[5883] = 8'h8;
        my_rom[5884] = 8'h8;
        my_rom[5885] = 8'h8;
        my_rom[5886] = 8'h8;
        my_rom[5887] = 8'h8;
        my_rom[5888] = 8'h8;
        my_rom[5889] = 8'h8;
        my_rom[5890] = 8'h8;
        my_rom[5891] = 8'ha;
        my_rom[5892] = 8'h8;
        my_rom[5893] = 8'h8;
        my_rom[5894] = 8'h8;
        my_rom[5895] = 8'h8;
        my_rom[5896] = 8'h8;
        my_rom[5897] = 8'h8;
        my_rom[5898] = 8'h8;
        my_rom[5899] = 8'h8;
        my_rom[5900] = 8'h8;
        my_rom[5901] = 8'h8;
        my_rom[5902] = 8'h8;
        my_rom[5903] = 8'h8;
        my_rom[5904] = 8'hf7;
        my_rom[5905] = 8'hf7;
        my_rom[5906] = 8'hf7;
        my_rom[5907] = 8'hf7;
        my_rom[5908] = 8'hed;
        my_rom[5909] = 8'had;
        my_rom[5910] = 8'had;
        my_rom[5911] = 8'hed;
        my_rom[5912] = 8'hed;
        my_rom[5913] = 8'hed;
        my_rom[5914] = 8'hed;
        my_rom[5915] = 8'hed;
        my_rom[5916] = 8'hed;
        my_rom[5917] = 8'hed;
        my_rom[5918] = 8'hef;
        my_rom[5919] = 8'hed;
        my_rom[5920] = 8'hef;
        my_rom[5921] = 8'hed;
        my_rom[5922] = 8'hed;
        my_rom[5923] = 8'hed;
        my_rom[5924] = 8'hed;
        my_rom[5925] = 8'ha5;
        my_rom[5926] = 8'ha5;
        my_rom[5927] = 8'ha5;
        my_rom[5928] = 8'ha5;
        my_rom[5929] = 8'ha5;
        my_rom[5930] = 8'ha5;
        my_rom[5931] = 8'ha5;
        my_rom[5932] = 8'ha5;
        my_rom[5933] = 8'ha5;
        my_rom[5934] = 8'ha5;
        my_rom[5935] = 8'ha5;
        my_rom[5936] = 8'ha5;
        my_rom[5937] = 8'h5b;
        my_rom[5938] = 8'h8;
        my_rom[5939] = 8'h8;
        my_rom[5940] = 8'h8;
        my_rom[5941] = 8'h8;
        my_rom[5942] = 8'h8;
        my_rom[5943] = 8'h8;
        my_rom[5944] = 8'h8;
        my_rom[5945] = 8'h8;
        my_rom[5946] = 8'h8;
        my_rom[5947] = 8'h8;
        my_rom[5948] = 8'h8;
        my_rom[5949] = 8'h8;
        my_rom[5950] = 8'h8;
        my_rom[5951] = 8'ha;
        my_rom[5952] = 8'h8;
        my_rom[5953] = 8'h8;
        my_rom[5954] = 8'h8;
        my_rom[5955] = 8'h8;
        my_rom[5956] = 8'h8;
        my_rom[5957] = 8'h8;
        my_rom[5958] = 8'h8;
        my_rom[5959] = 8'h8;
        my_rom[5960] = 8'h8;
        my_rom[5961] = 8'h8;
        my_rom[5962] = 8'h8;
        my_rom[5963] = 8'h8;
        my_rom[5964] = 8'h8;
        my_rom[5965] = 8'hf7;
        my_rom[5966] = 8'hf7;
        my_rom[5967] = 8'hf7;
        my_rom[5968] = 8'hf7;
        my_rom[5969] = 8'hed;
        my_rom[5970] = 8'had;
        my_rom[5971] = 8'had;
        my_rom[5972] = 8'had;
        my_rom[5973] = 8'hed;
        my_rom[5974] = 8'hed;
        my_rom[5975] = 8'hed;
        my_rom[5976] = 8'hed;
        my_rom[5977] = 8'hed;
        my_rom[5978] = 8'hed;
        my_rom[5979] = 8'hef;
        my_rom[5980] = 8'hef;
        my_rom[5981] = 8'hed;
        my_rom[5982] = 8'hed;
        my_rom[5983] = 8'hed;
        my_rom[5984] = 8'hed;
        my_rom[5985] = 8'ha5;
        my_rom[5986] = 8'ha5;
        my_rom[5987] = 8'ha5;
        my_rom[5988] = 8'ha5;
        my_rom[5989] = 8'ha5;
        my_rom[5990] = 8'ha5;
        my_rom[5991] = 8'ha5;
        my_rom[5992] = 8'had;
        my_rom[5993] = 8'ha5;
        my_rom[5994] = 8'ha5;
        my_rom[5995] = 8'ha5;
        my_rom[5996] = 8'h5b;
        my_rom[5997] = 8'h53;
        my_rom[5998] = 8'h8;
        my_rom[5999] = 8'h8;
        my_rom[6000] = 8'h8;
        my_rom[6001] = 8'h8;
        my_rom[6002] = 8'h8;
        my_rom[6003] = 8'h8;
        my_rom[6004] = 8'h8;
        my_rom[6005] = 8'h8;
        my_rom[6006] = 8'h8;
        my_rom[6007] = 8'h8;
        my_rom[6008] = 8'h8;
        my_rom[6009] = 8'h8;
        my_rom[6010] = 8'h8;
        my_rom[6011] = 8'ha;
        my_rom[6012] = 8'h8;
        my_rom[6013] = 8'h8;
        my_rom[6014] = 8'h8;
        my_rom[6015] = 8'h8;
        my_rom[6016] = 8'h8;
        my_rom[6017] = 8'h8;
        my_rom[6018] = 8'h8;
        my_rom[6019] = 8'h8;
        my_rom[6020] = 8'h8;
        my_rom[6021] = 8'h8;
        my_rom[6022] = 8'h8;
        my_rom[6023] = 8'h8;
        my_rom[6024] = 8'h8;
        my_rom[6025] = 8'h8;
        my_rom[6026] = 8'hf7;
        my_rom[6027] = 8'hf7;
        my_rom[6028] = 8'hf7;
        my_rom[6029] = 8'hf5;
        my_rom[6030] = 8'hed;
        my_rom[6031] = 8'had;
        my_rom[6032] = 8'ha5;
        my_rom[6033] = 8'had;
        my_rom[6034] = 8'had;
        my_rom[6035] = 8'hed;
        my_rom[6036] = 8'hed;
        my_rom[6037] = 8'hed;
        my_rom[6038] = 8'hed;
        my_rom[6039] = 8'hed;
        my_rom[6040] = 8'hed;
        my_rom[6041] = 8'hed;
        my_rom[6042] = 8'hed;
        my_rom[6043] = 8'ha5;
        my_rom[6044] = 8'ha5;
        my_rom[6045] = 8'ha5;
        my_rom[6046] = 8'ha5;
        my_rom[6047] = 8'ha5;
        my_rom[6048] = 8'ha5;
        my_rom[6049] = 8'ha5;
        my_rom[6050] = 8'ha5;
        my_rom[6051] = 8'ha5;
        my_rom[6052] = 8'ha5;
        my_rom[6053] = 8'ha5;
        my_rom[6054] = 8'ha5;
        my_rom[6055] = 8'ha3;
        my_rom[6056] = 8'h53;
        my_rom[6057] = 8'h8;
        my_rom[6058] = 8'h8;
        my_rom[6059] = 8'h8;
        my_rom[6060] = 8'h8;
        my_rom[6061] = 8'h8;
        my_rom[6062] = 8'h8;
        my_rom[6063] = 8'h8;
        my_rom[6064] = 8'h8;
        my_rom[6065] = 8'h8;
        my_rom[6066] = 8'h8;
        my_rom[6067] = 8'h8;
        my_rom[6068] = 8'h8;
        my_rom[6069] = 8'h8;
        my_rom[6070] = 8'h8;
        my_rom[6071] = 8'ha;
        my_rom[6072] = 8'h8;
        my_rom[6073] = 8'h8;
        my_rom[6074] = 8'h8;
        my_rom[6075] = 8'h8;
        my_rom[6076] = 8'h8;
        my_rom[6077] = 8'h8;
        my_rom[6078] = 8'h8;
        my_rom[6079] = 8'h8;
        my_rom[6080] = 8'h8;
        my_rom[6081] = 8'h8;
        my_rom[6082] = 8'h8;
        my_rom[6083] = 8'h8;
        my_rom[6084] = 8'h8;
        my_rom[6085] = 8'h8;
        my_rom[6086] = 8'h8;
        my_rom[6087] = 8'hf7;
        my_rom[6088] = 8'hf7;
        my_rom[6089] = 8'hf7;
        my_rom[6090] = 8'hf5;
        my_rom[6091] = 8'hed;
        my_rom[6092] = 8'had;
        my_rom[6093] = 8'ha5;
        my_rom[6094] = 8'ha5;
        my_rom[6095] = 8'ha5;
        my_rom[6096] = 8'had;
        my_rom[6097] = 8'had;
        my_rom[6098] = 8'had;
        my_rom[6099] = 8'had;
        my_rom[6100] = 8'ha5;
        my_rom[6101] = 8'ha5;
        my_rom[6102] = 8'ha5;
        my_rom[6103] = 8'ha5;
        my_rom[6104] = 8'h9b;
        my_rom[6105] = 8'h9b;
        my_rom[6106] = 8'h9b;
        my_rom[6107] = 8'h9b;
        my_rom[6108] = 8'h9b;
        my_rom[6109] = 8'ha3;
        my_rom[6110] = 8'ha3;
        my_rom[6111] = 8'ha5;
        my_rom[6112] = 8'ha5;
        my_rom[6113] = 8'ha5;
        my_rom[6114] = 8'had;
        my_rom[6115] = 8'ha5;
        my_rom[6116] = 8'h8;
        my_rom[6117] = 8'h8;
        my_rom[6118] = 8'h8;
        my_rom[6119] = 8'h8;
        my_rom[6120] = 8'h8;
        my_rom[6121] = 8'h8;
        my_rom[6122] = 8'h8;
        my_rom[6123] = 8'h8;
        my_rom[6124] = 8'h8;
        my_rom[6125] = 8'h8;
        my_rom[6126] = 8'h8;
        my_rom[6127] = 8'h8;
        my_rom[6128] = 8'h8;
        my_rom[6129] = 8'h8;
        my_rom[6130] = 8'h8;
        my_rom[6131] = 8'ha;
        my_rom[6132] = 8'h8;
        my_rom[6133] = 8'h8;
        my_rom[6134] = 8'h8;
        my_rom[6135] = 8'h8;
        my_rom[6136] = 8'h8;
        my_rom[6137] = 8'h8;
        my_rom[6138] = 8'h8;
        my_rom[6139] = 8'h8;
        my_rom[6140] = 8'h8;
        my_rom[6141] = 8'h8;
        my_rom[6142] = 8'h8;
        my_rom[6143] = 8'h8;
        my_rom[6144] = 8'h8;
        my_rom[6145] = 8'h8;
        my_rom[6146] = 8'h8;
        my_rom[6147] = 8'h8;
        my_rom[6148] = 8'hf7;
        my_rom[6149] = 8'hf7;
        my_rom[6150] = 8'hf5;
        my_rom[6151] = 8'hed;
        my_rom[6152] = 8'hed;
        my_rom[6153] = 8'had;
        my_rom[6154] = 8'ha5;
        my_rom[6155] = 8'ha5;
        my_rom[6156] = 8'ha5;
        my_rom[6157] = 8'ha5;
        my_rom[6158] = 8'ha5;
        my_rom[6159] = 8'ha5;
        my_rom[6160] = 8'ha5;
        my_rom[6161] = 8'ha3;
        my_rom[6162] = 8'h9b;
        my_rom[6163] = 8'h9b;
        my_rom[6164] = 8'h9b;
        my_rom[6165] = 8'h9b;
        my_rom[6166] = 8'h9b;
        my_rom[6167] = 8'h9b;
        my_rom[6168] = 8'h9b;
        my_rom[6169] = 8'h9b;
        my_rom[6170] = 8'h9b;
        my_rom[6171] = 8'h9b;
        my_rom[6172] = 8'ha3;
        my_rom[6173] = 8'had;
        my_rom[6174] = 8'had;
        my_rom[6175] = 8'h5b;
        my_rom[6176] = 8'h8;
        my_rom[6177] = 8'h8;
        my_rom[6178] = 8'h8;
        my_rom[6179] = 8'h8;
        my_rom[6180] = 8'h8;
        my_rom[6181] = 8'h8;
        my_rom[6182] = 8'h8;
        my_rom[6183] = 8'h8;
        my_rom[6184] = 8'h8;
        my_rom[6185] = 8'h8;
        my_rom[6186] = 8'h8;
        my_rom[6187] = 8'h8;
        my_rom[6188] = 8'h8;
        my_rom[6189] = 8'h8;
        my_rom[6190] = 8'h8;
        my_rom[6191] = 8'ha;
        my_rom[6192] = 8'h8;
        my_rom[6193] = 8'h8;
        my_rom[6194] = 8'h8;
        my_rom[6195] = 8'h8;
        my_rom[6196] = 8'h8;
        my_rom[6197] = 8'h8;
        my_rom[6198] = 8'h8;
        my_rom[6199] = 8'h8;
        my_rom[6200] = 8'h8;
        my_rom[6201] = 8'h8;
        my_rom[6202] = 8'h8;
        my_rom[6203] = 8'h8;
        my_rom[6204] = 8'h8;
        my_rom[6205] = 8'h8;
        my_rom[6206] = 8'h8;
        my_rom[6207] = 8'h8;
        my_rom[6208] = 8'h8;
        my_rom[6209] = 8'hf7;
        my_rom[6210] = 8'hf5;
        my_rom[6211] = 8'hf5;
        my_rom[6212] = 8'hed;
        my_rom[6213] = 8'hed;
        my_rom[6214] = 8'had;
        my_rom[6215] = 8'ha5;
        my_rom[6216] = 8'ha5;
        my_rom[6217] = 8'ha5;
        my_rom[6218] = 8'ha5;
        my_rom[6219] = 8'ha5;
        my_rom[6220] = 8'h9b;
        my_rom[6221] = 8'h9b;
        my_rom[6222] = 8'h9b;
        my_rom[6223] = 8'h9b;
        my_rom[6224] = 8'h9b;
        my_rom[6225] = 8'h93;
        my_rom[6226] = 8'h93;
        my_rom[6227] = 8'h93;
        my_rom[6228] = 8'h93;
        my_rom[6229] = 8'h9b;
        my_rom[6230] = 8'h9b;
        my_rom[6231] = 8'ha5;
        my_rom[6232] = 8'had;
        my_rom[6233] = 8'had;
        my_rom[6234] = 8'ha5;
        my_rom[6235] = 8'h5b;
        my_rom[6236] = 8'h8;
        my_rom[6237] = 8'h8;
        my_rom[6238] = 8'h8;
        my_rom[6239] = 8'h8;
        my_rom[6240] = 8'h8;
        my_rom[6241] = 8'h8;
        my_rom[6242] = 8'h8;
        my_rom[6243] = 8'h8;
        my_rom[6244] = 8'h8;
        my_rom[6245] = 8'h8;
        my_rom[6246] = 8'h8;
        my_rom[6247] = 8'h8;
        my_rom[6248] = 8'h8;
        my_rom[6249] = 8'h8;
        my_rom[6250] = 8'h8;
        my_rom[6251] = 8'ha;
        my_rom[6252] = 8'h8;
        my_rom[6253] = 8'h8;
        my_rom[6254] = 8'h8;
        my_rom[6255] = 8'h8;
        my_rom[6256] = 8'h8;
        my_rom[6257] = 8'h8;
        my_rom[6258] = 8'h8;
        my_rom[6259] = 8'h8;
        my_rom[6260] = 8'h8;
        my_rom[6261] = 8'h8;
        my_rom[6262] = 8'h8;
        my_rom[6263] = 8'h8;
        my_rom[6264] = 8'h8;
        my_rom[6265] = 8'h8;
        my_rom[6266] = 8'h8;
        my_rom[6267] = 8'h8;
        my_rom[6268] = 8'h8;
        my_rom[6269] = 8'h8;
        my_rom[6270] = 8'hf7;
        my_rom[6271] = 8'hf5;
        my_rom[6272] = 8'hf5;
        my_rom[6273] = 8'hed;
        my_rom[6274] = 8'hed;
        my_rom[6275] = 8'hed;
        my_rom[6276] = 8'ha5;
        my_rom[6277] = 8'ha3;
        my_rom[6278] = 8'h9b;
        my_rom[6279] = 8'h9b;
        my_rom[6280] = 8'h9b;
        my_rom[6281] = 8'h9b;
        my_rom[6282] = 8'h9b;
        my_rom[6283] = 8'h9b;
        my_rom[6284] = 8'h93;
        my_rom[6285] = 8'h93;
        my_rom[6286] = 8'h93;
        my_rom[6287] = 8'h93;
        my_rom[6288] = 8'h9b;
        my_rom[6289] = 8'h9b;
        my_rom[6290] = 8'ha5;
        my_rom[6291] = 8'ha5;
        my_rom[6292] = 8'had;
        my_rom[6293] = 8'had;
        my_rom[6294] = 8'haf;
        my_rom[6295] = 8'h8;
        my_rom[6296] = 8'h8;
        my_rom[6297] = 8'h8;
        my_rom[6298] = 8'h8;
        my_rom[6299] = 8'h8;
        my_rom[6300] = 8'h8;
        my_rom[6301] = 8'h8;
        my_rom[6302] = 8'h8;
        my_rom[6303] = 8'h8;
        my_rom[6304] = 8'h8;
        my_rom[6305] = 8'h8;
        my_rom[6306] = 8'h8;
        my_rom[6307] = 8'h8;
        my_rom[6308] = 8'h8;
        my_rom[6309] = 8'h8;
        my_rom[6310] = 8'h8;
        my_rom[6311] = 8'ha;
        my_rom[6312] = 8'h8;
        my_rom[6313] = 8'h8;
        my_rom[6314] = 8'h8;
        my_rom[6315] = 8'h8;
        my_rom[6316] = 8'h8;
        my_rom[6317] = 8'h8;
        my_rom[6318] = 8'h8;
        my_rom[6319] = 8'h8;
        my_rom[6320] = 8'h8;
        my_rom[6321] = 8'h8;
        my_rom[6322] = 8'h8;
        my_rom[6323] = 8'h8;
        my_rom[6324] = 8'h8;
        my_rom[6325] = 8'h8;
        my_rom[6326] = 8'h8;
        my_rom[6327] = 8'h8;
        my_rom[6328] = 8'h8;
        my_rom[6329] = 8'h8;
        my_rom[6330] = 8'h8;
        my_rom[6331] = 8'hf5;
        my_rom[6332] = 8'hf5;
        my_rom[6333] = 8'hed;
        my_rom[6334] = 8'hed;
        my_rom[6335] = 8'hed;
        my_rom[6336] = 8'had;
        my_rom[6337] = 8'ha5;
        my_rom[6338] = 8'ha3;
        my_rom[6339] = 8'h9b;
        my_rom[6340] = 8'h9b;
        my_rom[6341] = 8'h9b;
        my_rom[6342] = 8'h9b;
        my_rom[6343] = 8'h9b;
        my_rom[6344] = 8'h9b;
        my_rom[6345] = 8'h9b;
        my_rom[6346] = 8'h9b;
        my_rom[6347] = 8'h9b;
        my_rom[6348] = 8'h9b;
        my_rom[6349] = 8'ha5;
        my_rom[6350] = 8'ha5;
        my_rom[6351] = 8'had;
        my_rom[6352] = 8'had;
        my_rom[6353] = 8'had;
        my_rom[6354] = 8'haf;
        my_rom[6355] = 8'h8;
        my_rom[6356] = 8'h8;
        my_rom[6357] = 8'h8;
        my_rom[6358] = 8'h8;
        my_rom[6359] = 8'h8;
        my_rom[6360] = 8'h8;
        my_rom[6361] = 8'h8;
        my_rom[6362] = 8'h8;
        my_rom[6363] = 8'h8;
        my_rom[6364] = 8'h8;
        my_rom[6365] = 8'h8;
        my_rom[6366] = 8'h8;
        my_rom[6367] = 8'h8;
        my_rom[6368] = 8'h8;
        my_rom[6369] = 8'h8;
        my_rom[6370] = 8'h8;
        my_rom[6371] = 8'ha;
        my_rom[6372] = 8'h8;
        my_rom[6373] = 8'h8;
        my_rom[6374] = 8'h8;
        my_rom[6375] = 8'h8;
        my_rom[6376] = 8'h8;
        my_rom[6377] = 8'h8;
        my_rom[6378] = 8'h8;
        my_rom[6379] = 8'h8;
        my_rom[6380] = 8'h8;
        my_rom[6381] = 8'h8;
        my_rom[6382] = 8'h8;
        my_rom[6383] = 8'h8;
        my_rom[6384] = 8'h8;
        my_rom[6385] = 8'h8;
        my_rom[6386] = 8'h8;
        my_rom[6387] = 8'h8;
        my_rom[6388] = 8'h8;
        my_rom[6389] = 8'h8;
        my_rom[6390] = 8'h8;
        my_rom[6391] = 8'h8;
        my_rom[6392] = 8'hed;
        my_rom[6393] = 8'hed;
        my_rom[6394] = 8'hed;
        my_rom[6395] = 8'hed;
        my_rom[6396] = 8'hed;
        my_rom[6397] = 8'ha5;
        my_rom[6398] = 8'ha5;
        my_rom[6399] = 8'ha3;
        my_rom[6400] = 8'ha3;
        my_rom[6401] = 8'h9b;
        my_rom[6402] = 8'h9b;
        my_rom[6403] = 8'h9b;
        my_rom[6404] = 8'h9b;
        my_rom[6405] = 8'h9b;
        my_rom[6406] = 8'h9b;
        my_rom[6407] = 8'h9b;
        my_rom[6408] = 8'ha3;
        my_rom[6409] = 8'ha5;
        my_rom[6410] = 8'ha5;
        my_rom[6411] = 8'had;
        my_rom[6412] = 8'had;
        my_rom[6413] = 8'had;
        my_rom[6414] = 8'had;
        my_rom[6415] = 8'h8;
        my_rom[6416] = 8'h8;
        my_rom[6417] = 8'h8;
        my_rom[6418] = 8'h8;
        my_rom[6419] = 8'h8;
        my_rom[6420] = 8'h8;
        my_rom[6421] = 8'h8;
        my_rom[6422] = 8'h8;
        my_rom[6423] = 8'h8;
        my_rom[6424] = 8'h8;
        my_rom[6425] = 8'h8;
        my_rom[6426] = 8'h8;
        my_rom[6427] = 8'h8;
        my_rom[6428] = 8'h8;
        my_rom[6429] = 8'h8;
        my_rom[6430] = 8'h8;
        my_rom[6431] = 8'ha;
        my_rom[6432] = 8'h8;
        my_rom[6433] = 8'h8;
        my_rom[6434] = 8'h8;
        my_rom[6435] = 8'h8;
        my_rom[6436] = 8'h8;
        my_rom[6437] = 8'h8;
        my_rom[6438] = 8'h8;
        my_rom[6439] = 8'h8;
        my_rom[6440] = 8'h8;
        my_rom[6441] = 8'h8;
        my_rom[6442] = 8'h8;
        my_rom[6443] = 8'h8;
        my_rom[6444] = 8'h8;
        my_rom[6445] = 8'h8;
        my_rom[6446] = 8'h8;
        my_rom[6447] = 8'h8;
        my_rom[6448] = 8'h8;
        my_rom[6449] = 8'h8;
        my_rom[6450] = 8'h8;
        my_rom[6451] = 8'h8;
        my_rom[6452] = 8'h8;
        my_rom[6453] = 8'hed;
        my_rom[6454] = 8'hed;
        my_rom[6455] = 8'hed;
        my_rom[6456] = 8'hed;
        my_rom[6457] = 8'had;
        my_rom[6458] = 8'ha5;
        my_rom[6459] = 8'ha5;
        my_rom[6460] = 8'ha3;
        my_rom[6461] = 8'ha3;
        my_rom[6462] = 8'h9b;
        my_rom[6463] = 8'h9b;
        my_rom[6464] = 8'h9b;
        my_rom[6465] = 8'h9b;
        my_rom[6466] = 8'h9b;
        my_rom[6467] = 8'ha3;
        my_rom[6468] = 8'ha5;
        my_rom[6469] = 8'ha5;
        my_rom[6470] = 8'ha5;
        my_rom[6471] = 8'had;
        my_rom[6472] = 8'had;
        my_rom[6473] = 8'had;
        my_rom[6474] = 8'ha5;
        my_rom[6475] = 8'h8;
        my_rom[6476] = 8'h8;
        my_rom[6477] = 8'h8;
        my_rom[6478] = 8'h8;
        my_rom[6479] = 8'h8;
        my_rom[6480] = 8'h8;
        my_rom[6481] = 8'h8;
        my_rom[6482] = 8'h8;
        my_rom[6483] = 8'h8;
        my_rom[6484] = 8'h8;
        my_rom[6485] = 8'h8;
        my_rom[6486] = 8'h8;
        my_rom[6487] = 8'h8;
        my_rom[6488] = 8'h8;
        my_rom[6489] = 8'h8;
        my_rom[6490] = 8'h8;
        my_rom[6491] = 8'ha;
        my_rom[6492] = 8'h8;
        my_rom[6493] = 8'h8;
        my_rom[6494] = 8'h8;
        my_rom[6495] = 8'h8;
        my_rom[6496] = 8'h8;
        my_rom[6497] = 8'h8;
        my_rom[6498] = 8'h8;
        my_rom[6499] = 8'h8;
        my_rom[6500] = 8'h8;
        my_rom[6501] = 8'h8;
        my_rom[6502] = 8'h8;
        my_rom[6503] = 8'h8;
        my_rom[6504] = 8'h8;
        my_rom[6505] = 8'h8;
        my_rom[6506] = 8'h8;
        my_rom[6507] = 8'h8;
        my_rom[6508] = 8'h8;
        my_rom[6509] = 8'h8;
        my_rom[6510] = 8'h8;
        my_rom[6511] = 8'h8;
        my_rom[6512] = 8'h8;
        my_rom[6513] = 8'h8;
        my_rom[6514] = 8'h8;
        my_rom[6515] = 8'h8;
        my_rom[6516] = 8'h8;
        my_rom[6517] = 8'h8;
        my_rom[6518] = 8'h8;
        my_rom[6519] = 8'h8;
        my_rom[6520] = 8'h8;
        my_rom[6521] = 8'h8;
        my_rom[6522] = 8'h8;
        my_rom[6523] = 8'h8;
        my_rom[6524] = 8'h8;
        my_rom[6525] = 8'h8;
        my_rom[6526] = 8'h8;
        my_rom[6527] = 8'ha5;
        my_rom[6528] = 8'ha5;
        my_rom[6529] = 8'ha5;
        my_rom[6530] = 8'ha5;
        my_rom[6531] = 8'had;
        my_rom[6532] = 8'had;
        my_rom[6533] = 8'had;
        my_rom[6534] = 8'h5d;
        my_rom[6535] = 8'h8;
        my_rom[6536] = 8'h8;
        my_rom[6537] = 8'h8;
        my_rom[6538] = 8'h8;
        my_rom[6539] = 8'h8;
        my_rom[6540] = 8'h8;
        my_rom[6541] = 8'h8;
        my_rom[6542] = 8'h8;
        my_rom[6543] = 8'h8;
        my_rom[6544] = 8'h8;
        my_rom[6545] = 8'h8;
        my_rom[6546] = 8'h8;
        my_rom[6547] = 8'h8;
        my_rom[6548] = 8'h8;
        my_rom[6549] = 8'h8;
        my_rom[6550] = 8'h8;
        my_rom[6551] = 8'ha;
        my_rom[6552] = 8'hc;
    end
endmodule
